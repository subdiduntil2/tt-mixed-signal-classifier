magic
tech sky130A
magscale 1 2
timestamp 1755204415
<< viali >>
rect 2540 132 2578 172
rect 1600 64 1658 116
rect 2064 -854 2102 -818
<< metal1 >>
rect 1974 1296 2174 1496
rect 2034 1230 2128 1296
rect 1770 1182 2400 1230
rect 1772 732 1810 1182
rect 1988 900 2188 1100
rect 1772 714 1920 732
rect 1786 698 1920 714
rect 1690 416 1700 510
rect 1774 416 1784 510
rect 1936 436 1946 498
rect 2002 484 2012 498
rect 2054 484 2094 900
rect 2358 740 2400 1182
rect 2252 712 2400 740
rect 2252 706 2386 712
rect 2138 484 2148 508
rect 2002 452 2148 484
rect 2002 436 2012 452
rect 2138 440 2148 452
rect 2228 440 2238 508
rect 2398 436 2408 502
rect 2462 436 2472 502
rect 1810 300 1820 382
rect 1896 300 1906 382
rect 2052 310 2062 384
rect 2116 310 2126 384
rect 2280 294 2290 372
rect 2344 294 2354 372
rect 2610 286 2620 370
rect 2672 352 2682 370
rect 2752 352 2952 460
rect 2672 318 2952 352
rect 2672 312 2692 318
rect 2672 286 2682 312
rect 2752 260 2952 318
rect 2526 186 2568 188
rect 2526 172 3482 186
rect 2526 132 2540 172
rect 2578 158 3482 172
rect 2578 132 3476 158
rect 1632 128 1672 130
rect 548 116 1672 128
rect 548 64 1600 116
rect 1658 64 1672 116
rect 2526 112 3476 132
rect 2528 110 3476 112
rect 1784 76 1918 110
rect 2244 76 2378 110
rect 3370 84 3476 110
rect 548 48 1672 64
rect 556 -1126 668 48
rect 1632 46 1672 48
rect 1772 -130 1932 -96
rect 2260 -130 2394 -96
rect 910 -228 1110 -206
rect 910 -232 1212 -228
rect 910 -340 1130 -232
rect 1220 -340 1230 -232
rect 910 -406 1110 -340
rect 1806 -342 1816 -274
rect 1892 -342 1902 -274
rect 1670 -486 1680 -396
rect 1778 -486 1788 -396
rect 1922 -458 1932 -386
rect 1998 -396 2008 -386
rect 2050 -396 2060 -362
rect 1998 -458 2060 -396
rect 2050 -460 2060 -458
rect 2120 -396 2130 -362
rect 2120 -458 2198 -396
rect 2258 -410 2268 -280
rect 2368 -410 2378 -280
rect 2952 -402 2962 -310
rect 3024 -344 3034 -310
rect 3074 -344 3274 -206
rect 3024 -384 3274 -344
rect 3024 -402 3034 -384
rect 3074 -406 3274 -384
rect 2120 -460 2130 -458
rect 2160 -560 2170 -488
rect 2236 -560 2246 -488
rect 2394 -558 2404 -474
rect 2460 -558 2470 -474
rect 872 -726 1072 -612
rect 872 -728 1074 -726
rect 1766 -728 1926 -722
rect 872 -756 1926 -728
rect 2254 -730 2388 -726
rect 3036 -730 3236 -606
rect 872 -812 1072 -756
rect 2054 -818 2112 -738
rect 2254 -758 3236 -730
rect 2254 -760 2388 -758
rect 3036 -806 3236 -758
rect 2054 -854 2064 -818
rect 2102 -854 2112 -818
rect 2054 -1068 2112 -854
rect 2000 -1118 2200 -1068
rect 3370 -1112 3480 84
rect 3340 -1118 3480 -1112
rect 2000 -1126 3480 -1118
rect 204 -1190 3480 -1126
rect 2000 -1222 3480 -1190
rect 2000 -1226 3476 -1222
rect 2000 -1268 2200 -1226
<< via1 >>
rect 1700 416 1774 510
rect 1946 436 2002 498
rect 2148 440 2228 508
rect 2408 436 2462 502
rect 1820 300 1896 382
rect 2062 310 2116 384
rect 2290 294 2344 372
rect 2620 286 2672 370
rect 1130 -340 1220 -232
rect 1816 -342 1892 -274
rect 1680 -486 1778 -396
rect 1932 -458 1998 -386
rect 2060 -460 2120 -362
rect 2268 -410 2368 -280
rect 2962 -402 3024 -310
rect 2170 -560 2236 -488
rect 2404 -558 2460 -474
<< metal2 >>
rect 1700 510 1774 520
rect 2148 508 2228 518
rect 1946 498 2002 508
rect 1774 444 1946 486
rect 1946 426 2002 436
rect 2408 502 2462 512
rect 2228 452 2408 484
rect 2148 430 2228 440
rect 2408 426 2462 436
rect 1700 406 1774 416
rect 1820 382 1896 392
rect 2062 384 2116 394
rect 1896 318 2062 364
rect 1820 290 1896 300
rect 2060 310 2062 318
rect 1130 -232 1220 -222
rect 1816 -274 1892 -264
rect 1220 -324 1816 -282
rect 1130 -350 1220 -340
rect 1816 -352 1892 -342
rect 2060 -352 2116 310
rect 2290 372 2344 382
rect 2620 370 2672 380
rect 2344 302 2620 350
rect 2290 284 2344 294
rect 2620 276 2672 286
rect 2268 -280 2368 -270
rect 2060 -362 2120 -352
rect 1932 -386 1998 -376
rect 1680 -394 1778 -386
rect 1680 -396 1932 -394
rect 1778 -450 1932 -396
rect 1998 -446 2016 -394
rect 1932 -468 1998 -458
rect 2962 -310 3024 -300
rect 2368 -396 2962 -314
rect 2268 -420 2368 -410
rect 2962 -412 3024 -402
rect 2060 -470 2120 -460
rect 2404 -474 2460 -464
rect 1680 -496 1778 -486
rect 2170 -488 2236 -478
rect 2236 -542 2404 -498
rect 2170 -570 2236 -560
rect 2404 -568 2460 -558
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM1
timestamp 1754378775
transform 1 0 2315 0 1 407
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM3
timestamp 1754378775
transform 1 0 1851 0 1 -425
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM5
timestamp 1754378775
transform 1 0 2315 0 1 -425
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM8
timestamp 1754378775
transform 1 0 1851 0 1 407
box -285 -469 285 469
<< labels >>
flabel metal1 872 -812 1072 -612 0 FreeSans 256 0 0 0 Vin
port 4 nsew
flabel metal1 3036 -806 3236 -606 0 FreeSans 256 0 0 0 Vindot
port 5 nsew
flabel metal1 2752 260 2952 460 0 FreeSans 256 0 0 0 Vupper_out
port 1 nsew
flabel metal1 1988 900 2188 1100 0 FreeSans 256 0 0 0 Vupper
port 0 nsew
flabel metal1 1974 1296 2174 1496 0 FreeSans 256 0 0 0 Vg
port 2 nsew
flabel metal1 910 -406 1110 -206 0 FreeSans 256 0 0 0 Vout1
port 6 nsew
flabel metal1 3074 -406 3274 -206 0 FreeSans 256 0 0 0 Vout2
port 7 nsew
flabel metal1 2000 -1268 2200 -1068 0 FreeSans 256 0 0 0 Vdd
port 3 nsew
rlabel metal2 2070 28 2108 58 1 lmid
<< end >>
