VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_subdiduntil2_mixed_signal_classifier
  CLASS BLOCK ;
  FOREIGN tt_um_subdiduntil2_mixed_signal_classifier ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN VDPWR
    ANTENNAGATEAREA 3.006000 ;
    ANTENNADIFFAREA 124.248398 ;
    PORT
      LAYER nwell ;
        RECT 73.010 204.560 75.970 209.930 ;
        RECT 77.480 207.960 79.940 210.650 ;
        RECT 93.910 201.690 104.280 213.260 ;
        RECT 45.790 164.450 49.230 181.460 ;
        RECT 66.450 175.090 71.620 183.940 ;
        RECT 88.870 174.410 94.040 183.260 ;
        RECT 108.650 174.740 113.820 183.590 ;
        RECT 127.680 177.900 130.530 182.590 ;
        RECT 57.150 167.880 59.610 172.070 ;
        RECT 75.660 167.270 78.120 171.460 ;
        RECT 98.130 167.800 100.590 171.990 ;
        RECT 126.340 171.920 131.510 176.610 ;
        RECT 139.400 174.540 142.250 179.230 ;
        RECT 66.120 162.000 68.580 166.190 ;
        RECT 88.650 162.780 91.110 166.970 ;
        RECT 109.590 163.270 112.050 167.460 ;
        RECT 127.020 162.940 129.480 167.130 ;
        RECT 139.850 161.800 142.700 166.490 ;
        RECT 113.710 154.820 116.170 159.010 ;
        RECT 63.530 109.790 70.120 112.480 ;
        RECT 77.580 109.990 84.170 112.680 ;
        RECT 96.250 110.030 102.840 112.720 ;
        RECT 110.300 110.230 116.890 112.920 ;
        RECT 70.090 105.000 76.680 107.790 ;
        RECT 102.810 105.240 109.400 108.030 ;
        RECT 63.250 81.410 69.840 84.100 ;
        RECT 77.300 81.610 83.890 84.300 ;
        RECT 94.900 83.930 101.490 86.620 ;
        RECT 108.950 84.130 115.540 86.820 ;
        RECT 69.810 76.620 76.400 79.410 ;
        RECT 101.460 79.140 108.050 81.930 ;
        RECT 79.770 39.180 86.360 44.030 ;
      LAYER li1 ;
        RECT 91.570 214.300 103.950 214.840 ;
        RECT 98.050 213.080 98.270 213.130 ;
        RECT 101.400 213.080 101.580 213.170 ;
        RECT 94.090 212.910 104.100 213.080 ;
        RECT 77.950 210.470 78.170 210.510 ;
        RECT 77.660 210.300 79.760 210.470 ;
        RECT 75.240 209.750 75.440 209.840 ;
        RECT 73.190 209.580 75.790 209.750 ;
        RECT 73.190 204.910 73.360 209.580 ;
        RECT 75.050 207.815 75.220 208.855 ;
        RECT 75.050 205.635 75.220 206.675 ;
        RECT 75.620 204.910 75.790 209.580 ;
        RECT 77.660 208.310 77.830 210.300 ;
        RECT 78.230 209.035 78.400 209.575 ;
        RECT 79.590 208.310 79.760 210.300 ;
        RECT 77.660 208.140 79.760 208.310 ;
        RECT 94.090 209.400 94.260 212.910 ;
        RECT 96.550 211.725 96.720 212.185 ;
        RECT 96.550 210.125 96.720 210.585 ;
        RECT 99.010 209.400 99.180 212.910 ;
        RECT 103.930 209.400 104.100 212.910 ;
        RECT 94.090 209.230 104.100 209.400 ;
        RECT 94.090 208.940 94.300 209.230 ;
        RECT 94.090 205.840 94.260 208.940 ;
        RECT 94.020 205.720 94.260 205.840 ;
        RECT 99.010 205.720 99.180 209.230 ;
        RECT 103.930 205.720 104.100 209.230 ;
        RECT 94.020 205.550 104.100 205.720 ;
        RECT 94.020 205.460 94.260 205.550 ;
        RECT 73.190 204.740 75.790 204.910 ;
        RECT 94.090 202.040 94.260 205.460 ;
        RECT 99.010 202.040 99.180 205.550 ;
        RECT 103.930 202.040 104.100 205.550 ;
        RECT 94.090 201.870 104.100 202.040 ;
        RECT 66.630 183.590 71.440 183.760 ;
        RECT 45.970 181.110 49.050 181.280 ;
        RECT 45.970 164.800 46.140 181.110 ;
        RECT 47.130 179.925 47.300 180.385 ;
        RECT 48.310 179.925 48.480 180.385 ;
        RECT 47.130 178.325 47.300 178.785 ;
        RECT 48.310 178.325 48.480 178.785 ;
        RECT 47.130 176.725 47.300 177.185 ;
        RECT 48.310 176.725 48.480 177.185 ;
        RECT 47.130 175.125 47.300 175.585 ;
        RECT 48.310 175.125 48.480 175.585 ;
        RECT 48.880 174.060 49.050 181.110 ;
        RECT 66.630 180.140 66.800 183.590 ;
        RECT 67.200 180.325 67.370 182.865 ;
        RECT 68.380 180.325 68.550 182.865 ;
        RECT 66.620 179.880 66.910 180.140 ;
        RECT 66.630 179.600 66.800 179.880 ;
        RECT 68.950 179.600 69.120 183.590 ;
        RECT 69.520 180.325 69.690 182.865 ;
        RECT 70.700 180.325 70.870 182.865 ;
        RECT 71.270 180.420 71.440 183.590 ;
        RECT 108.830 183.240 113.640 183.410 ;
        RECT 89.050 182.910 93.860 183.080 ;
        RECT 71.270 180.220 71.510 180.420 ;
        RECT 71.270 179.600 71.440 180.220 ;
        RECT 66.630 179.430 71.440 179.600 ;
        RECT 89.050 179.460 89.220 182.910 ;
        RECT 66.630 175.440 66.800 179.430 ;
        RECT 68.950 175.470 69.120 179.430 ;
        RECT 68.940 175.440 69.130 175.470 ;
        RECT 71.270 175.440 71.440 179.430 ;
        RECT 89.040 179.200 89.330 179.460 ;
        RECT 66.630 175.270 71.440 175.440 ;
        RECT 89.050 178.920 89.220 179.200 ;
        RECT 91.370 178.920 91.540 182.910 ;
        RECT 93.690 179.740 93.860 182.910 ;
        RECT 108.830 179.790 109.000 183.240 ;
        RECT 93.690 179.540 93.930 179.740 ;
        RECT 93.690 178.920 93.860 179.540 ;
        RECT 108.820 179.530 109.110 179.790 ;
        RECT 89.050 178.750 93.860 178.920 ;
        RECT 89.050 174.760 89.220 178.750 ;
        RECT 91.370 174.790 91.540 178.750 ;
        RECT 91.360 174.760 91.550 174.790 ;
        RECT 93.690 174.760 93.860 178.750 ;
        RECT 108.830 179.250 109.000 179.530 ;
        RECT 111.150 179.250 111.320 183.240 ;
        RECT 113.470 180.070 113.640 183.240 ;
        RECT 126.650 182.920 131.840 183.320 ;
        RECT 129.140 182.410 129.330 182.450 ;
        RECT 127.860 182.240 130.350 182.410 ;
        RECT 113.470 179.870 113.710 180.070 ;
        RECT 113.470 179.250 113.640 179.870 ;
        RECT 108.830 179.080 113.640 179.250 ;
        RECT 108.830 175.090 109.000 179.080 ;
        RECT 111.150 175.120 111.320 179.080 ;
        RECT 111.140 175.090 111.330 175.120 ;
        RECT 113.470 175.090 113.640 179.080 ;
        RECT 127.860 178.250 128.030 182.240 ;
        RECT 130.180 178.250 130.350 182.240 ;
        RECT 139.550 179.050 139.760 179.080 ;
        RECT 139.550 178.880 142.070 179.050 ;
        RECT 139.550 178.700 139.760 178.880 ;
        RECT 127.860 178.080 130.350 178.250 ;
        RECT 127.000 176.430 127.180 176.480 ;
        RECT 130.960 176.430 131.170 176.510 ;
        RECT 108.830 174.920 113.640 175.090 ;
        RECT 126.520 176.260 131.330 176.430 ;
        RECT 89.050 174.590 93.860 174.760 ;
        RECT 48.880 174.050 49.170 174.060 ;
        RECT 47.130 173.525 47.300 173.985 ;
        RECT 48.310 173.525 48.480 173.985 ;
        RECT 48.820 173.320 49.170 174.050 ;
        RECT 47.130 171.925 47.300 172.385 ;
        RECT 48.310 171.925 48.480 172.385 ;
        RECT 47.130 170.325 47.300 170.785 ;
        RECT 48.310 170.325 48.480 170.785 ;
        RECT 47.130 168.725 47.300 169.185 ;
        RECT 48.310 168.725 48.480 169.185 ;
        RECT 47.130 167.125 47.300 167.585 ;
        RECT 48.310 167.125 48.480 167.585 ;
        RECT 47.130 165.525 47.300 165.985 ;
        RECT 48.310 165.525 48.480 165.985 ;
        RECT 48.880 164.800 49.050 173.320 ;
        RECT 126.520 172.270 126.690 176.260 ;
        RECT 128.840 172.270 129.010 176.260 ;
        RECT 131.160 172.270 131.330 176.260 ;
        RECT 139.580 174.890 139.750 178.700 ;
        RECT 141.900 174.890 142.070 178.880 ;
        RECT 139.580 174.720 142.070 174.890 ;
        RECT 126.520 172.100 131.330 172.270 ;
        RECT 57.330 171.720 59.430 171.890 ;
        RECT 57.330 169.990 57.500 171.720 ;
        RECT 57.330 169.650 57.570 169.990 ;
        RECT 57.330 168.230 57.500 169.650 ;
        RECT 57.900 168.955 58.070 170.995 ;
        RECT 59.260 168.230 59.430 171.720 ;
        RECT 98.310 171.640 100.410 171.810 ;
        RECT 57.330 168.060 59.430 168.230 ;
        RECT 75.840 171.110 77.940 171.280 ;
        RECT 75.840 169.380 76.010 171.110 ;
        RECT 75.840 169.040 76.080 169.380 ;
        RECT 75.840 167.620 76.010 169.040 ;
        RECT 76.410 168.345 76.580 170.385 ;
        RECT 77.770 167.620 77.940 171.110 ;
        RECT 98.310 169.910 98.480 171.640 ;
        RECT 98.310 169.570 98.550 169.910 ;
        RECT 98.310 168.150 98.480 169.570 ;
        RECT 98.880 168.875 99.050 170.915 ;
        RECT 100.240 168.150 100.410 171.640 ;
        RECT 98.310 167.980 100.410 168.150 ;
        RECT 75.840 167.450 77.940 167.620 ;
        RECT 109.770 167.110 111.870 167.280 ;
        RECT 88.830 166.620 90.930 166.790 ;
        RECT 45.970 164.630 49.050 164.800 ;
        RECT 66.300 165.840 68.400 166.010 ;
        RECT 66.300 164.110 66.470 165.840 ;
        RECT 66.300 163.770 66.540 164.110 ;
        RECT 66.300 162.350 66.470 163.770 ;
        RECT 66.870 163.075 67.040 165.115 ;
        RECT 68.230 162.350 68.400 165.840 ;
        RECT 88.830 164.890 89.000 166.620 ;
        RECT 88.830 164.550 89.070 164.890 ;
        RECT 88.830 163.130 89.000 164.550 ;
        RECT 89.400 163.855 89.570 165.895 ;
        RECT 90.760 163.130 90.930 166.620 ;
        RECT 109.770 165.380 109.940 167.110 ;
        RECT 109.770 165.040 110.010 165.380 ;
        RECT 109.770 163.620 109.940 165.040 ;
        RECT 110.340 164.345 110.510 166.385 ;
        RECT 111.700 163.620 111.870 167.110 ;
        RECT 109.770 163.450 111.870 163.620 ;
        RECT 127.200 166.780 129.300 166.950 ;
        RECT 127.200 165.050 127.370 166.780 ;
        RECT 127.200 164.710 127.440 165.050 ;
        RECT 88.830 162.960 90.930 163.130 ;
        RECT 127.200 163.290 127.370 164.710 ;
        RECT 127.770 164.015 127.940 166.055 ;
        RECT 129.130 163.290 129.300 166.780 ;
        RECT 140.030 166.140 142.520 166.310 ;
        RECT 140.030 165.970 140.200 166.140 ;
        RECT 139.990 165.700 140.200 165.970 ;
        RECT 127.200 163.120 129.300 163.290 ;
        RECT 66.300 162.180 68.400 162.350 ;
        RECT 140.030 162.150 140.200 165.700 ;
        RECT 142.350 162.150 142.520 166.140 ;
        RECT 140.030 161.980 142.520 162.150 ;
        RECT 46.815 160.320 47.145 160.490 ;
        RECT 47.405 160.320 47.735 160.490 ;
        RECT 47.995 160.320 48.325 160.490 ;
        RECT 113.890 158.660 115.990 158.830 ;
        RECT 46.815 158.100 47.145 158.270 ;
        RECT 47.405 158.100 47.735 158.270 ;
        RECT 47.995 158.100 48.325 158.270 ;
        RECT 46.815 157.560 47.145 157.730 ;
        RECT 47.405 157.560 47.735 157.730 ;
        RECT 47.995 157.560 48.325 157.730 ;
        RECT 113.890 156.930 114.060 158.660 ;
        RECT 113.890 156.590 114.130 156.930 ;
        RECT 46.815 155.340 47.145 155.510 ;
        RECT 47.405 155.340 47.735 155.510 ;
        RECT 47.995 155.340 48.325 155.510 ;
        RECT 113.890 155.170 114.060 156.590 ;
        RECT 114.460 155.895 114.630 157.935 ;
        RECT 115.820 155.170 115.990 158.660 ;
        RECT 113.890 155.000 115.990 155.170 ;
        RECT 64.970 113.840 80.560 114.560 ;
        RECT 97.690 114.080 113.280 114.800 ;
        RECT 113.500 112.740 113.710 112.780 ;
        RECT 110.480 112.570 116.710 112.740 ;
        RECT 99.460 112.540 99.630 112.550 ;
        RECT 80.780 112.500 80.990 112.540 ;
        RECT 77.760 112.330 83.990 112.500 ;
        RECT 66.740 112.300 66.910 112.310 ;
        RECT 63.710 112.130 69.940 112.300 ;
        RECT 63.710 110.140 63.880 112.130 ;
        RECT 66.170 110.865 66.340 111.405 ;
        RECT 66.740 110.140 66.910 112.130 ;
        RECT 67.310 110.865 67.480 111.405 ;
        RECT 69.770 110.140 69.940 112.130 ;
        RECT 77.760 110.340 77.930 112.330 ;
        RECT 80.220 111.065 80.390 111.605 ;
        RECT 80.790 110.340 80.960 112.330 ;
        RECT 81.360 111.065 81.530 111.605 ;
        RECT 83.820 110.340 83.990 112.330 ;
        RECT 77.760 110.170 83.990 110.340 ;
        RECT 96.430 112.370 102.660 112.540 ;
        RECT 96.430 110.380 96.600 112.370 ;
        RECT 98.890 111.105 99.060 111.645 ;
        RECT 99.460 110.380 99.630 112.370 ;
        RECT 100.030 111.105 100.200 111.645 ;
        RECT 102.490 110.380 102.660 112.370 ;
        RECT 110.480 110.580 110.650 112.570 ;
        RECT 112.940 111.305 113.110 111.845 ;
        RECT 113.510 110.580 113.680 112.570 ;
        RECT 114.080 111.305 114.250 111.845 ;
        RECT 116.540 110.580 116.710 112.570 ;
        RECT 110.480 110.410 116.710 110.580 ;
        RECT 96.430 110.210 102.660 110.380 ;
        RECT 63.710 109.970 69.940 110.140 ;
        RECT 106.000 107.850 106.270 107.900 ;
        RECT 102.990 107.680 109.220 107.850 ;
        RECT 73.280 107.610 73.550 107.660 ;
        RECT 70.270 107.440 76.500 107.610 ;
        RECT 70.270 105.350 70.440 107.440 ;
        RECT 73.300 105.350 73.470 107.440 ;
        RECT 76.330 105.350 76.500 107.440 ;
        RECT 102.990 105.590 103.160 107.680 ;
        RECT 106.020 105.590 106.190 107.680 ;
        RECT 109.050 105.590 109.220 107.680 ;
        RECT 102.990 105.420 109.220 105.590 ;
        RECT 70.270 105.180 76.500 105.350 ;
        RECT 96.340 87.980 111.930 88.700 ;
        RECT 112.150 86.640 112.360 86.680 ;
        RECT 109.130 86.470 115.360 86.640 ;
        RECT 98.110 86.440 98.280 86.450 ;
        RECT 95.080 86.270 101.310 86.440 ;
        RECT 64.690 85.460 80.280 86.180 ;
        RECT 95.080 84.280 95.250 86.270 ;
        RECT 97.540 85.005 97.710 85.545 ;
        RECT 98.110 84.280 98.280 86.270 ;
        RECT 98.680 85.005 98.850 85.545 ;
        RECT 101.140 84.280 101.310 86.270 ;
        RECT 109.130 84.480 109.300 86.470 ;
        RECT 111.590 85.205 111.760 85.745 ;
        RECT 112.160 84.480 112.330 86.470 ;
        RECT 112.730 85.205 112.900 85.745 ;
        RECT 115.190 84.480 115.360 86.470 ;
        RECT 109.130 84.310 115.360 84.480 ;
        RECT 80.500 84.120 80.710 84.160 ;
        RECT 77.480 83.950 83.710 84.120 ;
        RECT 95.080 84.110 101.310 84.280 ;
        RECT 66.460 83.920 66.630 83.930 ;
        RECT 63.430 83.750 69.660 83.920 ;
        RECT 63.430 81.760 63.600 83.750 ;
        RECT 65.890 82.485 66.060 83.025 ;
        RECT 66.460 81.760 66.630 83.750 ;
        RECT 67.030 82.485 67.200 83.025 ;
        RECT 69.490 81.760 69.660 83.750 ;
        RECT 77.480 81.960 77.650 83.950 ;
        RECT 79.940 82.685 80.110 83.225 ;
        RECT 80.510 81.960 80.680 83.950 ;
        RECT 81.080 82.685 81.250 83.225 ;
        RECT 83.540 81.960 83.710 83.950 ;
        RECT 77.480 81.790 83.710 81.960 ;
        RECT 63.430 81.590 69.660 81.760 ;
        RECT 104.650 81.750 104.920 81.800 ;
        RECT 101.640 81.580 107.870 81.750 ;
        RECT 101.640 79.490 101.810 81.580 ;
        RECT 104.670 79.490 104.840 81.580 ;
        RECT 107.700 79.490 107.870 81.580 ;
        RECT 101.640 79.320 107.870 79.490 ;
        RECT 73.000 79.230 73.270 79.280 ;
        RECT 69.990 79.060 76.220 79.230 ;
        RECT 69.990 76.970 70.160 79.060 ;
        RECT 73.020 76.970 73.190 79.060 ;
        RECT 76.050 76.970 76.220 79.060 ;
        RECT 69.990 76.800 76.220 76.970 ;
        RECT 82.920 43.850 83.240 43.910 ;
        RECT 79.950 43.680 86.180 43.850 ;
        RECT 79.950 41.690 80.120 43.680 ;
        RECT 82.410 42.415 82.580 42.955 ;
        RECT 82.980 41.710 83.150 43.680 ;
        RECT 83.550 42.415 83.720 42.955 ;
        RECT 82.940 41.690 83.200 41.710 ;
        RECT 86.010 41.690 86.180 43.680 ;
        RECT 79.950 41.520 86.180 41.690 ;
        RECT 79.950 39.530 80.120 41.520 ;
        RECT 82.980 39.530 83.150 41.520 ;
        RECT 86.010 39.530 86.180 41.520 ;
        RECT 79.950 39.360 86.180 39.530 ;
      LAYER met1 ;
        RECT 90.920 214.840 91.920 215.050 ;
        RECT 90.920 214.760 103.950 214.840 ;
        RECT 89.170 214.720 103.950 214.760 ;
        RECT 89.170 214.530 103.960 214.720 ;
        RECT 89.140 214.420 103.960 214.530 ;
        RECT 89.140 214.360 103.950 214.420 ;
        RECT 73.650 212.090 74.650 212.390 ;
        RECT 89.140 212.220 89.820 214.360 ;
        RECT 90.920 214.300 103.950 214.360 ;
        RECT 90.920 214.050 91.920 214.300 ;
        RECT 93.520 213.670 93.890 214.300 ;
        RECT 96.380 214.060 96.940 214.300 ;
        RECT 75.120 212.090 75.520 212.120 ;
        RECT 79.170 212.090 89.820 212.220 ;
        RECT 73.650 211.650 89.820 212.090 ;
        RECT 73.650 211.390 74.650 211.650 ;
        RECT 75.120 210.180 75.520 211.650 ;
        RECT 75.150 208.835 75.510 210.180 ;
        RECT 77.890 209.555 78.300 211.650 ;
        RECT 79.170 211.600 89.820 211.650 ;
        RECT 89.140 211.570 89.820 211.600 ;
        RECT 93.490 209.560 93.890 213.670 ;
        RECT 96.320 213.620 97.030 214.060 ;
        RECT 97.950 213.310 98.380 214.300 ;
        RECT 97.920 213.250 98.380 213.310 ;
        RECT 97.920 213.000 98.410 213.250 ;
        RECT 97.930 212.940 98.410 213.000 ;
        RECT 97.930 212.920 98.390 212.940 ;
        RECT 101.360 212.920 101.610 214.300 ;
        RECT 96.520 212.150 96.750 212.165 ;
        RECT 96.450 211.770 96.830 212.150 ;
        RECT 96.520 211.745 96.750 211.770 ;
        RECT 96.470 210.200 96.840 210.600 ;
        RECT 96.520 210.145 96.750 210.200 ;
        RECT 77.890 209.130 78.430 209.555 ;
        RECT 78.200 209.055 78.430 209.130 ;
        RECT 75.020 207.835 75.510 208.835 ;
        RECT 93.490 208.900 94.430 209.560 ;
        RECT 93.490 208.720 93.860 208.900 ;
        RECT 94.240 208.890 94.430 208.900 ;
        RECT 93.470 208.450 93.870 208.720 ;
        RECT 75.150 206.655 75.510 207.835 ;
        RECT 75.020 205.830 75.510 206.655 ;
        RECT 93.460 205.960 93.880 208.450 ;
        RECT 75.020 205.655 75.250 205.830 ;
        RECT 93.440 205.360 94.430 205.960 ;
        RECT 46.590 187.420 49.820 190.060 ;
        RECT 48.460 185.840 48.990 187.420 ;
        RECT 48.470 184.830 48.990 185.840 ;
        RECT 55.500 184.830 56.180 184.920 ;
        RECT 48.470 184.170 56.180 184.830 ;
        RECT 48.470 183.830 48.990 184.170 ;
        RECT 55.500 184.130 56.180 184.170 ;
        RECT 68.560 184.060 69.560 185.060 ;
        RECT 48.460 182.280 48.990 183.830 ;
        RECT 48.470 180.400 48.990 182.280 ;
        RECT 67.170 182.110 67.400 182.845 ;
        RECT 67.070 181.640 67.540 182.110 ;
        RECT 68.350 182.050 68.580 182.845 ;
        RECT 68.300 181.980 68.680 182.050 ;
        RECT 68.890 181.980 69.090 184.060 ;
        RECT 125.960 183.320 126.960 183.420 ;
        RECT 125.960 183.200 131.840 183.320 ;
        RECT 125.960 183.190 132.240 183.200 ;
        RECT 125.960 183.060 132.640 183.190 ;
        RECT 124.330 183.040 132.640 183.060 ;
        RECT 124.330 182.920 131.840 183.040 ;
        RECT 69.490 182.100 69.720 182.845 ;
        RECT 69.310 181.980 69.810 182.100 ;
        RECT 70.670 182.070 70.900 182.845 ;
        RECT 124.330 182.670 126.960 182.920 ;
        RECT 68.300 181.820 69.810 181.980 ;
        RECT 68.300 181.740 68.680 181.820 ;
        RECT 69.310 181.760 69.810 181.820 ;
        RECT 48.440 180.370 48.990 180.400 ;
        RECT 48.290 180.365 48.990 180.370 ;
        RECT 47.100 180.330 47.330 180.365 ;
        RECT 47.000 180.000 47.370 180.330 ;
        RECT 47.100 179.945 47.330 180.000 ;
        RECT 48.280 179.945 48.990 180.365 ;
        RECT 67.170 180.345 67.400 181.640 ;
        RECT 68.350 180.345 68.580 181.740 ;
        RECT 69.490 180.345 69.720 181.760 ;
        RECT 70.610 181.740 70.980 182.070 ;
        RECT 70.670 180.345 70.900 181.740 ;
        RECT 71.250 180.490 71.460 180.500 ;
        RECT 66.780 180.200 66.980 180.210 ;
        RECT 48.290 179.920 48.990 179.945 ;
        RECT 48.440 179.820 48.990 179.920 ;
        RECT 48.440 178.780 48.870 179.820 ;
        RECT 61.360 179.800 66.980 180.200 ;
        RECT 71.250 180.120 76.030 180.490 ;
        RECT 124.330 180.260 124.710 182.670 ;
        RECT 125.960 182.420 126.960 182.670 ;
        RECT 128.970 182.580 129.430 182.920 ;
        RECT 128.980 182.330 129.430 182.580 ;
        RECT 128.980 182.140 129.440 182.330 ;
        RECT 71.260 180.110 76.030 180.120 ;
        RECT 48.300 178.765 48.870 178.780 ;
        RECT 47.100 178.750 47.330 178.765 ;
        RECT 46.990 178.420 47.360 178.750 ;
        RECT 47.100 178.345 47.330 178.420 ;
        RECT 48.280 178.345 48.870 178.765 ;
        RECT 48.300 178.330 48.870 178.345 ;
        RECT 48.440 177.690 48.870 178.330 ;
        RECT 48.440 177.620 48.940 177.690 ;
        RECT 48.440 177.600 49.010 177.620 ;
        RECT 48.450 177.420 49.010 177.600 ;
        RECT 48.450 177.400 48.940 177.420 ;
        RECT 48.440 177.380 48.940 177.400 ;
        RECT 48.440 177.180 48.870 177.380 ;
        RECT 47.100 177.130 47.330 177.165 ;
        RECT 47.040 176.800 47.410 177.130 ;
        RECT 47.100 176.745 47.330 176.800 ;
        RECT 48.260 176.730 48.870 177.180 ;
        RECT 48.440 175.570 48.870 176.730 ;
        RECT 47.100 175.520 47.330 175.565 ;
        RECT 47.020 175.190 47.390 175.520 ;
        RECT 47.100 175.145 47.330 175.190 ;
        RECT 48.230 175.120 48.870 175.570 ;
        RECT 48.440 174.220 48.870 175.120 ;
        RECT 61.400 174.220 61.960 179.800 ;
        RECT 66.780 179.790 66.980 179.800 ;
        RECT 75.470 179.950 76.030 180.110 ;
        RECT 113.450 180.140 113.660 180.150 ;
        RECT 117.570 180.140 124.710 180.260 ;
        RECT 68.890 174.220 69.180 175.870 ;
        RECT 75.470 174.220 76.020 179.950 ;
        RECT 108.980 179.850 109.180 179.860 ;
        RECT 93.670 179.810 93.880 179.820 ;
        RECT 93.670 179.670 98.450 179.810 ;
        RECT 89.200 179.520 89.400 179.530 ;
        RECT 83.780 179.120 89.400 179.520 ;
        RECT 93.670 179.440 98.420 179.670 ;
        RECT 103.560 179.450 109.180 179.850 ;
        RECT 113.450 179.770 124.710 180.140 ;
        RECT 113.460 179.760 124.710 179.770 ;
        RECT 117.570 179.680 124.710 179.760 ;
        RECT 93.680 179.430 98.420 179.440 ;
        RECT 48.440 173.990 76.050 174.220 ;
        RECT 47.100 173.920 47.330 173.965 ;
        RECT 47.040 173.590 47.410 173.920 ;
        RECT 47.100 173.545 47.330 173.590 ;
        RECT 48.250 173.580 76.050 173.990 ;
        RECT 83.820 173.580 84.380 179.120 ;
        RECT 89.200 179.110 89.400 179.120 ;
        RECT 97.890 179.300 98.420 179.430 ;
        RECT 48.250 173.540 88.560 173.580 ;
        RECT 91.310 173.540 91.600 175.190 ;
        RECT 48.440 173.510 97.680 173.540 ;
        RECT 97.890 173.510 98.440 179.300 ;
        RECT 103.600 173.580 104.160 179.450 ;
        RECT 108.980 179.440 109.180 179.450 ;
        RECT 111.090 173.870 111.380 175.520 ;
        RECT 110.820 173.620 111.820 173.870 ;
        RECT 117.670 173.730 118.530 179.680 ;
        RECT 124.330 178.500 124.710 179.680 ;
        RECT 132.330 179.200 132.630 183.040 ;
        RECT 130.910 178.940 139.840 179.200 ;
        RECT 130.890 178.560 139.840 178.940 ;
        RECT 130.890 178.530 132.770 178.560 ;
        RECT 124.330 178.330 127.230 178.500 ;
        RECT 124.330 178.180 127.240 178.330 ;
        RECT 126.920 176.700 127.240 178.180 ;
        RECT 126.840 176.250 127.240 176.700 ;
        RECT 130.890 176.240 131.310 178.530 ;
        RECT 117.140 173.620 119.400 173.730 ;
        RECT 110.820 173.580 119.400 173.620 ;
        RECT 101.840 173.510 119.400 173.580 ;
        RECT 48.440 173.120 119.400 173.510 ;
        RECT 48.440 172.370 48.870 173.120 ;
        RECT 47.100 172.310 47.330 172.365 ;
        RECT 47.020 171.980 47.390 172.310 ;
        RECT 47.100 171.945 47.330 171.980 ;
        RECT 48.230 171.920 48.870 172.370 ;
        RECT 48.440 170.765 48.870 171.920 ;
        RECT 47.100 170.690 47.330 170.765 ;
        RECT 48.280 170.730 48.870 170.765 ;
        RECT 46.980 170.390 47.360 170.690 ;
        RECT 47.100 170.345 47.330 170.390 ;
        RECT 48.240 170.380 48.870 170.730 ;
        RECT 48.280 170.345 48.870 170.380 ;
        RECT 48.440 169.190 48.870 170.345 ;
        RECT 47.100 169.130 47.330 169.165 ;
        RECT 47.000 168.800 47.370 169.130 ;
        RECT 47.100 168.745 47.330 168.800 ;
        RECT 48.270 168.740 48.870 169.190 ;
        RECT 48.440 167.600 48.870 168.740 ;
        RECT 47.100 167.550 47.330 167.565 ;
        RECT 47.000 167.220 47.370 167.550 ;
        RECT 47.100 167.145 47.330 167.220 ;
        RECT 48.230 167.150 48.870 167.600 ;
        RECT 48.280 167.145 48.870 167.150 ;
        RECT 48.440 165.990 48.870 167.145 ;
        RECT 47.100 165.920 47.330 165.965 ;
        RECT 46.980 165.590 47.350 165.920 ;
        RECT 48.260 165.610 48.870 165.990 ;
        RECT 47.100 165.545 47.330 165.590 ;
        RECT 48.260 165.540 48.670 165.610 ;
        RECT 51.000 161.220 52.600 173.120 ;
        RECT 55.560 170.320 56.430 173.120 ;
        RECT 55.520 170.070 56.520 170.320 ;
        RECT 57.870 170.070 58.100 170.975 ;
        RECT 55.520 169.610 58.100 170.070 ;
        RECT 55.520 169.320 56.520 169.610 ;
        RECT 57.870 168.975 58.100 169.610 ;
        RECT 64.530 164.440 65.550 173.120 ;
        RECT 74.050 173.080 119.400 173.120 ;
        RECT 74.050 172.870 111.820 173.080 ;
        RECT 117.140 173.010 119.400 173.080 ;
        RECT 74.050 172.840 111.020 172.870 ;
        RECT 74.050 172.820 106.390 172.840 ;
        RECT 74.050 172.810 88.560 172.820 ;
        RECT 74.050 169.710 74.920 172.810 ;
        RECT 74.030 169.460 75.030 169.710 ;
        RECT 76.380 169.460 76.610 170.365 ;
        RECT 74.030 169.000 76.610 169.460 ;
        RECT 74.030 168.710 75.030 169.000 ;
        RECT 76.380 168.365 76.610 169.000 ;
        RECT 64.490 164.190 65.550 164.440 ;
        RECT 66.840 164.190 67.070 165.095 ;
        RECT 87.020 164.970 88.070 172.810 ;
        RECT 91.040 172.750 106.390 172.820 ;
        RECT 91.040 172.540 92.040 172.750 ;
        RECT 96.450 172.740 106.390 172.750 ;
        RECT 107.860 172.740 111.020 172.840 ;
        RECT 96.450 170.240 97.410 172.740 ;
        RECT 96.450 169.990 97.500 170.240 ;
        RECT 98.850 169.990 99.080 170.895 ;
        RECT 96.450 169.530 99.080 169.990 ;
        RECT 96.450 169.240 97.500 169.530 ;
        RECT 96.450 169.170 97.410 169.240 ;
        RECT 98.850 168.895 99.080 169.530 ;
        RECT 89.370 164.970 89.600 165.875 ;
        RECT 108.140 165.710 108.830 172.740 ;
        RECT 87.020 164.510 89.600 164.970 ;
        RECT 107.960 165.460 108.960 165.710 ;
        RECT 110.310 165.460 110.540 166.365 ;
        RECT 118.810 165.500 119.400 173.010 ;
        RECT 107.960 165.000 110.540 165.460 ;
        RECT 107.960 164.710 108.960 165.000 ;
        RECT 87.020 164.440 88.070 164.510 ;
        RECT 87.020 164.220 88.020 164.440 ;
        RECT 64.490 163.730 67.070 164.190 ;
        RECT 89.370 163.875 89.600 164.510 ;
        RECT 110.310 164.365 110.540 165.000 ;
        RECT 118.570 165.170 119.400 165.500 ;
        RECT 125.390 165.170 126.390 165.380 ;
        RECT 118.570 165.130 126.390 165.170 ;
        RECT 127.740 165.130 127.970 166.035 ;
        RECT 137.830 166.030 138.440 178.560 ;
        RECT 137.830 165.600 140.300 166.030 ;
        RECT 118.570 164.760 127.970 165.130 ;
        RECT 64.490 163.720 65.550 163.730 ;
        RECT 64.490 163.440 65.490 163.720 ;
        RECT 66.840 163.095 67.070 163.730 ;
        RECT 48.120 161.200 52.620 161.220 ;
        RECT 48.100 161.070 52.620 161.200 ;
        RECT 48.100 160.520 48.240 161.070 ;
        RECT 46.835 160.490 47.125 160.520 ;
        RECT 47.425 160.490 47.715 160.520 ;
        RECT 48.015 160.490 48.305 160.520 ;
        RECT 46.835 160.300 48.305 160.490 ;
        RECT 46.835 160.290 47.125 160.300 ;
        RECT 47.425 160.290 47.715 160.300 ;
        RECT 48.015 160.290 48.305 160.300 ;
        RECT 46.835 158.250 47.125 158.300 ;
        RECT 47.425 158.250 47.715 158.300 ;
        RECT 48.015 158.250 48.305 158.300 ;
        RECT 46.835 158.140 48.305 158.250 ;
        RECT 51.000 158.140 52.600 161.070 ;
        RECT 118.570 159.550 119.330 164.760 ;
        RECT 125.390 164.670 127.970 164.760 ;
        RECT 125.390 164.380 126.390 164.670 ;
        RECT 127.740 164.035 127.970 164.670 ;
        RECT 112.210 159.300 119.330 159.550 ;
        RECT 46.835 158.070 52.600 158.140 ;
        RECT 46.840 157.760 52.600 158.070 ;
        RECT 46.835 157.570 52.600 157.760 ;
        RECT 112.130 159.090 119.330 159.300 ;
        RECT 112.130 159.040 119.270 159.090 ;
        RECT 46.835 157.540 48.305 157.570 ;
        RECT 46.835 157.530 47.125 157.540 ;
        RECT 47.425 157.530 47.715 157.540 ;
        RECT 48.015 157.530 48.305 157.540 ;
        RECT 46.835 155.510 47.125 155.540 ;
        RECT 47.425 155.510 47.715 155.540 ;
        RECT 48.015 155.510 48.305 155.540 ;
        RECT 46.835 155.320 48.305 155.510 ;
        RECT 46.835 155.310 47.125 155.320 ;
        RECT 47.410 154.600 47.720 155.320 ;
        RECT 48.015 155.310 48.305 155.320 ;
        RECT 51.920 154.660 52.590 157.570 ;
        RECT 112.130 157.260 112.890 159.040 ;
        RECT 112.080 157.010 113.080 157.260 ;
        RECT 114.430 157.010 114.660 157.915 ;
        RECT 112.080 156.550 114.660 157.010 ;
        RECT 112.080 156.260 113.080 156.550 ;
        RECT 114.430 155.915 114.660 156.550 ;
        RECT 47.140 153.940 47.860 154.600 ;
        RECT 51.820 154.560 52.590 154.660 ;
        RECT 51.820 153.890 52.560 154.560 ;
        RECT 113.490 114.960 113.810 114.980 ;
        RECT 97.170 114.940 113.810 114.960 ;
        RECT 80.770 114.720 81.090 114.740 ;
        RECT 64.450 114.700 81.090 114.720 ;
        RECT 63.680 113.700 81.090 114.700 ;
        RECT 96.400 113.940 113.810 114.940 ;
        RECT 97.170 113.910 113.810 113.940 ;
        RECT 64.450 113.670 81.090 113.700 ;
        RECT 66.140 111.250 66.370 111.385 ;
        RECT 66.680 111.250 66.940 113.670 ;
        RECT 67.280 111.250 67.510 111.385 ;
        RECT 66.140 111.070 67.510 111.250 ;
        RECT 70.430 111.190 70.640 113.670 ;
        RECT 80.190 111.460 80.420 111.585 ;
        RECT 80.570 111.460 81.100 113.670 ;
        RECT 81.330 111.460 81.560 111.585 ;
        RECT 66.140 110.885 66.370 111.070 ;
        RECT 67.280 110.885 67.510 111.070 ;
        RECT 70.390 110.770 70.790 111.190 ;
        RECT 80.190 111.170 81.560 111.460 ;
        RECT 73.060 110.610 73.830 111.160 ;
        RECT 80.190 111.085 80.420 111.170 ;
        RECT 81.330 111.085 81.560 111.170 ;
        RECT 98.860 111.490 99.090 111.625 ;
        RECT 99.400 111.490 99.660 113.910 ;
        RECT 100.000 111.490 100.230 111.625 ;
        RECT 98.860 111.310 100.230 111.490 ;
        RECT 103.150 111.430 103.360 113.910 ;
        RECT 112.910 111.700 113.140 111.825 ;
        RECT 113.290 111.700 113.820 113.910 ;
        RECT 114.050 111.700 114.280 111.825 ;
        RECT 98.860 111.125 99.090 111.310 ;
        RECT 100.000 111.125 100.230 111.310 ;
        RECT 103.110 111.010 103.510 111.430 ;
        RECT 112.910 111.410 114.280 111.700 ;
        RECT 105.780 110.850 106.550 111.400 ;
        RECT 112.910 111.325 113.140 111.410 ;
        RECT 114.050 111.325 114.280 111.410 ;
        RECT 73.170 107.270 73.720 110.610 ;
        RECT 105.890 107.510 106.440 110.850 ;
        RECT 118.110 88.910 119.110 89.060 ;
        RECT 111.750 88.860 119.110 88.910 ;
        RECT 95.820 88.840 119.110 88.860 ;
        RECT 95.050 88.060 119.110 88.840 ;
        RECT 95.050 88.010 118.710 88.060 ;
        RECT 95.050 87.840 112.460 88.010 ;
        RECT 95.820 87.810 112.460 87.840 ;
        RECT 80.490 86.340 80.810 86.360 ;
        RECT 64.170 86.320 80.810 86.340 ;
        RECT 63.400 85.320 80.810 86.320 ;
        RECT 64.170 85.290 80.810 85.320 ;
        RECT 97.510 85.390 97.740 85.525 ;
        RECT 98.050 85.390 98.310 87.810 ;
        RECT 98.650 85.390 98.880 85.525 ;
        RECT 65.860 82.870 66.090 83.005 ;
        RECT 66.400 82.870 66.660 85.290 ;
        RECT 67.000 82.870 67.230 83.005 ;
        RECT 65.860 82.690 67.230 82.870 ;
        RECT 70.150 82.810 70.360 85.290 ;
        RECT 79.910 83.080 80.140 83.205 ;
        RECT 80.290 83.080 80.820 85.290 ;
        RECT 97.510 85.210 98.880 85.390 ;
        RECT 101.800 85.330 102.010 87.810 ;
        RECT 111.560 85.600 111.790 85.725 ;
        RECT 111.940 85.600 112.470 87.810 ;
        RECT 112.700 85.600 112.930 85.725 ;
        RECT 97.510 85.025 97.740 85.210 ;
        RECT 98.650 85.025 98.880 85.210 ;
        RECT 101.760 84.910 102.160 85.330 ;
        RECT 111.560 85.310 112.930 85.600 ;
        RECT 104.430 84.750 105.200 85.300 ;
        RECT 111.560 85.225 111.790 85.310 ;
        RECT 112.700 85.225 112.930 85.310 ;
        RECT 81.050 83.080 81.280 83.205 ;
        RECT 65.860 82.505 66.090 82.690 ;
        RECT 67.000 82.505 67.230 82.690 ;
        RECT 70.110 82.390 70.510 82.810 ;
        RECT 79.910 82.790 81.280 83.080 ;
        RECT 72.780 82.230 73.550 82.780 ;
        RECT 79.910 82.705 80.140 82.790 ;
        RECT 81.050 82.705 81.280 82.790 ;
        RECT 72.890 78.890 73.440 82.230 ;
        RECT 104.540 81.410 105.090 84.750 ;
        RECT 82.580 44.390 83.720 45.370 ;
        RECT 82.660 44.370 83.660 44.390 ;
        RECT 82.380 42.810 82.610 42.935 ;
        RECT 82.850 42.810 83.300 44.370 ;
        RECT 83.520 42.810 83.750 42.935 ;
        RECT 82.380 42.640 83.750 42.810 ;
        RECT 82.380 42.435 82.610 42.640 ;
        RECT 82.870 41.430 83.300 42.640 ;
        RECT 83.520 42.435 83.750 42.640 ;
      LAYER met2 ;
        RECT 90.980 214.070 91.760 215.000 ;
        RECT 96.370 213.570 96.980 214.110 ;
        RECT 96.560 212.200 96.870 213.570 ;
        RECT 96.500 211.920 96.870 212.200 ;
        RECT 96.500 211.720 96.780 211.920 ;
        RECT 96.570 210.650 96.710 211.720 ;
        RECT 96.520 210.150 96.790 210.650 ;
        RECT 46.640 187.370 49.770 190.110 ;
        RECT 55.550 184.730 56.130 184.970 ;
        RECT 68.680 184.730 69.470 184.860 ;
        RECT 55.550 184.130 69.490 184.730 ;
        RECT 55.550 184.080 56.130 184.130 ;
        RECT 67.120 181.990 67.490 182.160 ;
        RECT 68.350 181.990 68.630 182.100 ;
        RECT 67.120 181.780 68.630 181.990 ;
        RECT 67.120 181.590 67.490 181.780 ;
        RECT 68.350 181.690 68.630 181.780 ;
        RECT 69.360 181.980 69.760 182.150 ;
        RECT 70.660 181.980 70.930 182.120 ;
        RECT 69.360 181.820 70.930 181.980 ;
        RECT 69.360 181.710 69.760 181.820 ;
        RECT 70.660 181.690 70.930 181.820 ;
        RECT 47.000 179.800 47.450 180.490 ;
        RECT 48.240 179.810 48.690 180.500 ;
        RECT 46.940 178.220 47.390 178.910 ;
        RECT 48.250 178.240 48.700 178.930 ;
        RECT 46.970 176.640 47.420 177.330 ;
        RECT 48.240 176.640 48.690 177.330 ;
        RECT 47.030 175.010 47.480 175.700 ;
        RECT 48.220 175.010 48.670 175.700 ;
        RECT 46.970 173.430 47.420 174.120 ;
        RECT 48.240 173.410 48.690 174.100 ;
        RECT 46.980 171.810 47.410 172.480 ;
        RECT 48.220 171.820 48.650 172.490 ;
        RECT 46.980 170.270 47.470 170.860 ;
        RECT 48.190 170.280 48.670 170.870 ;
        RECT 46.990 168.630 47.440 169.320 ;
        RECT 48.210 168.650 48.660 169.340 ;
        RECT 46.970 167.020 47.420 167.710 ;
        RECT 48.200 167.010 48.650 167.700 ;
        RECT 46.930 165.420 47.380 166.110 ;
        RECT 48.240 165.410 48.690 166.100 ;
        RECT 47.190 154.520 47.810 154.650 ;
        RECT 51.870 154.520 52.510 154.710 ;
        RECT 47.190 153.970 52.560 154.520 ;
        RECT 47.190 153.890 47.810 153.970 ;
        RECT 51.870 153.840 52.510 153.970 ;
        RECT 64.630 113.690 65.390 114.720 ;
        RECT 97.570 113.860 98.300 114.720 ;
        RECT 103.160 111.390 103.460 111.480 ;
        RECT 105.830 111.390 106.500 111.450 ;
        RECT 70.440 111.150 70.740 111.240 ;
        RECT 73.110 111.150 73.780 111.210 ;
        RECT 70.440 110.790 73.780 111.150 ;
        RECT 103.160 111.030 106.500 111.390 ;
        RECT 103.160 110.960 103.460 111.030 ;
        RECT 105.830 110.800 106.500 111.030 ;
        RECT 70.440 110.720 70.740 110.790 ;
        RECT 73.110 110.560 73.780 110.790 ;
        RECT 95.680 87.930 96.420 88.740 ;
        RECT 65.200 85.390 66.160 86.300 ;
        RECT 101.810 85.290 102.110 85.380 ;
        RECT 104.480 85.290 105.150 85.350 ;
        RECT 101.810 84.930 105.150 85.290 ;
        RECT 101.810 84.860 102.110 84.930 ;
        RECT 104.480 84.700 105.150 84.930 ;
        RECT 70.160 82.770 70.460 82.860 ;
        RECT 72.830 82.770 73.500 82.830 ;
        RECT 70.160 82.410 73.500 82.770 ;
        RECT 70.160 82.340 70.460 82.410 ;
        RECT 72.830 82.180 73.500 82.410 ;
        RECT 82.630 44.340 83.670 45.420 ;
      LAYER met3 ;
        RECT 90.930 214.095 91.810 214.975 ;
        RECT 46.590 187.395 49.820 190.085 ;
        RECT 46.950 180.380 47.500 180.465 ;
        RECT 48.190 180.380 48.740 180.475 ;
        RECT 46.950 179.930 48.740 180.380 ;
        RECT 46.950 179.825 47.500 179.930 ;
        RECT 48.190 179.835 48.740 179.930 ;
        RECT 46.890 178.800 47.440 178.885 ;
        RECT 48.200 178.800 48.750 178.905 ;
        RECT 46.890 178.350 48.750 178.800 ;
        RECT 46.890 178.245 47.440 178.350 ;
        RECT 48.200 178.265 48.750 178.350 ;
        RECT 46.920 177.190 47.470 177.305 ;
        RECT 48.190 177.190 48.740 177.305 ;
        RECT 46.920 176.740 48.740 177.190 ;
        RECT 46.920 176.665 47.470 176.740 ;
        RECT 48.190 176.665 48.740 176.740 ;
        RECT 46.980 175.600 47.530 175.675 ;
        RECT 48.170 175.600 48.720 175.675 ;
        RECT 46.980 175.150 48.720 175.600 ;
        RECT 46.980 175.035 47.530 175.150 ;
        RECT 48.170 175.035 48.720 175.150 ;
        RECT 46.920 173.920 47.470 174.095 ;
        RECT 48.190 173.920 48.740 174.075 ;
        RECT 46.920 173.580 48.740 173.920 ;
        RECT 46.920 173.455 47.470 173.580 ;
        RECT 48.190 173.435 48.740 173.580 ;
        RECT 46.930 172.310 47.460 172.455 ;
        RECT 48.170 172.310 48.700 172.465 ;
        RECT 46.930 171.990 48.700 172.310 ;
        RECT 46.930 171.835 47.460 171.990 ;
        RECT 48.170 171.845 48.700 171.990 ;
        RECT 46.930 170.770 47.520 170.835 ;
        RECT 48.140 170.770 48.720 170.845 ;
        RECT 46.930 170.380 48.720 170.770 ;
        RECT 46.930 170.295 47.520 170.380 ;
        RECT 48.140 170.305 48.720 170.380 ;
        RECT 46.940 169.140 47.490 169.295 ;
        RECT 48.160 169.140 48.710 169.315 ;
        RECT 46.940 168.820 48.710 169.140 ;
        RECT 46.940 168.655 47.490 168.820 ;
        RECT 48.160 168.675 48.710 168.820 ;
        RECT 46.920 167.530 47.470 167.685 ;
        RECT 48.150 167.530 48.700 167.675 ;
        RECT 46.920 167.210 48.700 167.530 ;
        RECT 46.920 167.045 47.470 167.210 ;
        RECT 48.150 167.035 48.700 167.210 ;
        RECT 46.880 165.990 47.430 166.085 ;
        RECT 48.190 165.990 48.740 166.075 ;
        RECT 46.880 165.680 48.740 165.990 ;
        RECT 46.880 165.445 47.430 165.680 ;
        RECT 48.190 165.435 48.740 165.680 ;
        RECT 64.580 113.715 65.440 114.695 ;
        RECT 97.520 113.885 98.350 114.695 ;
        RECT 95.630 87.955 96.470 88.715 ;
        RECT 65.200 86.275 66.260 86.280 ;
        RECT 65.150 85.470 66.260 86.275 ;
        RECT 65.150 85.415 66.210 85.470 ;
        RECT 82.580 44.365 83.720 45.395 ;
      LAYER met4 ;
        RECT 26.510 214.880 28.510 219.730 ;
        RECT 31.460 214.880 34.990 214.970 ;
        RECT 26.510 214.850 36.970 214.880 ;
        RECT 50.030 214.850 57.760 214.910 ;
        RECT 90.975 214.850 91.765 214.955 ;
        RECT 26.510 213.850 95.620 214.850 ;
        RECT 26.510 213.660 36.970 213.850 ;
        RECT 50.030 213.830 57.760 213.850 ;
        RECT 26.510 191.380 28.510 213.660 ;
        RECT 31.460 213.590 34.990 213.660 ;
        RECT 26.510 189.580 28.390 191.380 ;
        RECT 46.635 189.580 49.775 190.065 ;
        RECT 26.510 189.490 50.010 189.580 ;
        RECT 26.410 187.540 50.010 189.490 ;
        RECT 26.410 187.500 28.390 187.540 ;
        RECT 26.510 187.090 28.390 187.500 ;
        RECT 46.635 187.415 49.775 187.540 ;
        RECT 26.510 170.540 28.510 187.090 ;
        RECT 26.510 168.590 28.280 170.540 ;
        RECT 26.510 114.800 28.510 168.590 ;
        RECT 31.460 114.800 35.550 115.100 ;
        RECT 26.510 114.540 35.550 114.800 ;
        RECT 64.625 114.540 65.395 114.675 ;
        RECT 97.565 114.540 98.305 114.675 ;
        RECT 26.510 113.980 98.790 114.540 ;
        RECT 26.510 113.780 65.840 113.980 ;
        RECT 97.565 113.905 98.305 113.980 ;
        RECT 26.510 113.490 35.550 113.780 ;
        RECT 64.625 113.735 65.395 113.780 ;
        RECT 26.510 87.240 28.510 113.490 ;
        RECT 31.460 113.210 35.550 113.490 ;
        RECT 64.920 88.050 99.930 88.860 ;
        RECT 26.370 86.460 38.590 87.240 ;
        RECT 65.090 86.460 66.320 88.050 ;
        RECT 95.675 87.975 96.425 88.050 ;
        RECT 26.370 85.170 66.590 86.460 ;
        RECT 26.370 84.540 38.590 85.170 ;
        RECT 26.510 46.130 28.510 84.540 ;
        RECT 26.510 45.450 40.080 46.130 ;
        RECT 26.510 43.840 85.380 45.450 ;
        RECT 26.510 43.430 40.080 43.840 ;
        RECT 26.510 3.970 28.510 43.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END VDPWR
  PIN VGND
    ANTENNAGATEAREA 2.688000 ;
    ANTENNADIFFAREA 39.495998 ;
    PORT
      LAYER pwell ;
        RECT 77.500 204.910 79.960 207.510 ;
        RECT 69.490 100.180 76.080 103.480 ;
        RECT 102.210 100.420 108.800 103.720 ;
        RECT 64.340 95.430 70.930 97.950 ;
        RECT 97.060 95.670 103.650 98.190 ;
        RECT 69.210 71.800 75.800 75.100 ;
        RECT 100.860 74.320 107.450 77.620 ;
        RECT 95.710 69.570 102.300 72.090 ;
        RECT 64.060 67.050 70.650 69.570 ;
        RECT 71.590 55.160 78.180 59.830 ;
        RECT 86.000 54.000 92.590 58.670 ;
      LAYER li1 ;
        RECT 77.680 207.160 79.780 207.330 ;
        RECT 77.680 205.260 77.850 207.160 ;
        RECT 78.250 205.940 78.420 206.480 ;
        RECT 78.060 205.260 78.280 205.380 ;
        RECT 79.610 205.260 79.780 207.160 ;
        RECT 77.680 205.090 79.780 205.260 ;
        RECT 99.810 205.040 101.410 205.210 ;
        RECT 101.700 205.040 103.300 205.210 ;
        RECT 101.470 204.365 101.640 204.825 ;
        RECT 99.810 203.980 101.410 204.150 ;
        RECT 101.700 203.980 103.300 204.150 ;
        RECT 99.810 203.440 101.410 203.610 ;
        RECT 101.700 203.440 103.300 203.610 ;
        RECT 101.470 202.765 101.640 203.225 ;
        RECT 99.810 202.380 101.410 202.550 ;
        RECT 101.700 202.380 103.300 202.550 ;
        RECT 92.770 200.430 104.690 200.950 ;
        RECT 102.390 103.370 108.620 103.540 ;
        RECT 69.670 103.130 75.900 103.300 ;
        RECT 69.670 100.530 69.840 103.130 ;
        RECT 72.700 100.550 72.870 103.130 ;
        RECT 72.670 100.530 72.900 100.550 ;
        RECT 75.730 100.530 75.900 103.130 ;
        RECT 102.390 100.770 102.560 103.370 ;
        RECT 105.420 100.790 105.590 103.370 ;
        RECT 105.390 100.770 105.620 100.790 ;
        RECT 108.450 100.770 108.620 103.370 ;
        RECT 102.390 100.600 108.620 100.770 ;
        RECT 69.670 100.360 75.900 100.530 ;
        RECT 97.240 97.840 103.470 98.010 ;
        RECT 64.520 97.600 70.750 97.770 ;
        RECT 64.520 95.780 64.690 97.600 ;
        RECT 66.980 96.460 67.150 96.920 ;
        RECT 67.550 95.830 67.720 97.600 ;
        RECT 68.120 96.460 68.290 96.920 ;
        RECT 67.550 95.780 67.740 95.830 ;
        RECT 70.580 95.780 70.750 97.600 ;
        RECT 97.240 96.020 97.410 97.840 ;
        RECT 99.700 96.700 99.870 97.160 ;
        RECT 100.270 96.070 100.440 97.840 ;
        RECT 100.840 96.700 101.010 97.160 ;
        RECT 100.270 96.020 100.460 96.070 ;
        RECT 103.300 96.020 103.470 97.840 ;
        RECT 97.240 95.850 103.470 96.020 ;
        RECT 64.520 95.610 70.750 95.780 ;
        RECT 64.460 93.590 85.330 93.850 ;
        RECT 97.180 93.830 118.050 94.090 ;
        RECT 101.040 77.270 107.270 77.440 ;
        RECT 69.390 74.750 75.620 74.920 ;
        RECT 69.390 72.150 69.560 74.750 ;
        RECT 72.420 72.170 72.590 74.750 ;
        RECT 72.390 72.150 72.620 72.170 ;
        RECT 75.450 72.150 75.620 74.750 ;
        RECT 101.040 74.670 101.210 77.270 ;
        RECT 104.070 74.690 104.240 77.270 ;
        RECT 104.040 74.670 104.270 74.690 ;
        RECT 107.100 74.670 107.270 77.270 ;
        RECT 101.040 74.500 107.270 74.670 ;
        RECT 69.390 71.980 75.620 72.150 ;
        RECT 95.890 71.740 102.120 71.910 ;
        RECT 95.890 69.920 96.060 71.740 ;
        RECT 98.350 70.600 98.520 71.060 ;
        RECT 98.920 69.970 99.090 71.740 ;
        RECT 99.490 70.600 99.660 71.060 ;
        RECT 98.920 69.920 99.110 69.970 ;
        RECT 101.950 69.920 102.120 71.740 ;
        RECT 95.890 69.750 102.120 69.920 ;
        RECT 64.240 69.220 70.470 69.390 ;
        RECT 64.240 67.400 64.410 69.220 ;
        RECT 66.700 68.080 66.870 68.540 ;
        RECT 67.270 67.450 67.440 69.220 ;
        RECT 67.840 68.080 68.010 68.540 ;
        RECT 67.270 67.400 67.460 67.450 ;
        RECT 70.300 67.400 70.470 69.220 ;
        RECT 95.830 67.730 116.700 67.990 ;
        RECT 64.240 67.230 70.470 67.400 ;
        RECT 64.180 65.210 85.050 65.470 ;
        RECT 71.770 59.480 78.000 59.650 ;
        RECT 71.770 57.580 71.940 59.480 ;
        RECT 74.800 57.600 74.970 59.480 ;
        RECT 74.800 57.580 75.010 57.600 ;
        RECT 77.830 57.580 78.000 59.480 ;
        RECT 71.770 57.410 78.000 57.580 ;
        RECT 71.770 55.510 71.940 57.410 ;
        RECT 74.230 56.190 74.400 56.730 ;
        RECT 74.800 55.560 74.970 57.410 ;
        RECT 75.370 56.190 75.540 56.730 ;
        RECT 74.800 55.510 75.100 55.560 ;
        RECT 77.830 55.510 78.000 57.410 ;
        RECT 71.770 55.340 78.000 55.510 ;
        RECT 86.180 58.320 92.410 58.490 ;
        RECT 86.180 56.420 86.350 58.320 ;
        RECT 89.210 56.440 89.380 58.320 ;
        RECT 89.210 56.420 89.420 56.440 ;
        RECT 92.240 56.420 92.410 58.320 ;
        RECT 86.180 56.250 92.410 56.420 ;
        RECT 74.810 55.330 75.100 55.340 ;
        RECT 86.180 54.350 86.350 56.250 ;
        RECT 88.640 55.030 88.810 55.570 ;
        RECT 89.210 54.400 89.380 56.250 ;
        RECT 89.780 55.030 89.950 55.570 ;
        RECT 89.210 54.350 89.510 54.400 ;
        RECT 92.240 54.350 92.410 56.250 ;
        RECT 86.180 54.180 92.410 54.350 ;
        RECT 89.220 54.170 89.510 54.180 ;
        RECT 78.710 19.850 88.550 21.665 ;
        RECT 90.480 19.920 100.320 21.735 ;
        RECT 78.630 19.680 88.630 19.850 ;
        RECT 90.400 19.750 100.400 19.920 ;
        RECT 77.330 17.060 89.660 17.780 ;
        RECT 90.680 17.010 100.580 17.760 ;
      LAYER met1 ;
        RECT 78.220 206.440 78.450 206.460 ;
        RECT 77.970 205.960 78.450 206.440 ;
        RECT 77.970 204.620 78.340 205.960 ;
        RECT 99.830 205.010 101.390 205.240 ;
        RECT 101.720 205.010 103.280 205.240 ;
        RECT 100.480 204.740 100.800 205.010 ;
        RECT 101.440 204.790 101.670 204.805 ;
        RECT 101.380 204.740 101.770 204.790 ;
        RECT 77.610 203.620 78.610 204.620 ;
        RECT 100.480 204.470 101.770 204.740 ;
        RECT 100.480 204.180 100.800 204.470 ;
        RECT 101.380 204.430 101.770 204.470 ;
        RECT 101.440 204.385 101.670 204.430 ;
        RECT 102.340 204.180 102.660 205.010 ;
        RECT 99.830 204.170 101.390 204.180 ;
        RECT 101.720 204.170 103.280 204.180 ;
        RECT 99.830 203.970 103.280 204.170 ;
        RECT 99.830 203.950 101.390 203.970 ;
        RECT 101.720 203.950 103.280 203.970 ;
        RECT 100.490 203.640 100.790 203.950 ;
        RECT 102.360 203.640 102.660 203.950 ;
        RECT 77.880 201.630 78.400 203.620 ;
        RECT 99.830 203.610 101.390 203.640 ;
        RECT 101.720 203.610 103.280 203.640 ;
        RECT 99.830 203.410 103.280 203.610 ;
        RECT 100.510 202.580 100.830 203.410 ;
        RECT 101.350 202.850 101.740 203.210 ;
        RECT 101.440 202.785 101.670 202.850 ;
        RECT 102.300 202.580 102.620 203.410 ;
        RECT 99.830 202.350 101.390 202.580 ;
        RECT 101.720 202.350 103.280 202.580 ;
        RECT 77.320 200.920 79.080 201.630 ;
        RECT 101.300 201.200 101.860 201.550 ;
        RECT 92.390 201.140 92.780 201.180 ;
        RECT 92.120 200.950 93.120 201.140 ;
        RECT 101.410 200.950 101.650 201.200 ;
        RECT 92.120 200.920 104.690 200.950 ;
        RECT 77.320 200.440 104.690 200.920 ;
        RECT 77.320 199.760 79.080 200.440 ;
        RECT 92.120 200.430 104.690 200.440 ;
        RECT 92.120 200.140 93.120 200.430 ;
        RECT 72.620 99.420 72.990 100.660 ;
        RECT 105.340 99.660 105.710 100.900 ;
        RECT 66.950 96.810 67.180 96.900 ;
        RECT 68.090 96.810 68.320 96.900 ;
        RECT 66.950 96.640 68.320 96.810 ;
        RECT 66.950 96.480 67.180 96.640 ;
        RECT 62.780 94.060 64.640 94.380 ;
        RECT 67.510 94.060 67.820 96.640 ;
        RECT 68.090 96.480 68.320 96.640 ;
        RECT 72.610 94.060 72.990 99.420 ;
        RECT 99.670 97.050 99.900 97.140 ;
        RECT 100.810 97.050 101.040 97.140 ;
        RECT 99.670 96.880 101.040 97.050 ;
        RECT 99.670 96.720 99.900 96.880 ;
        RECT 95.440 94.300 97.300 94.600 ;
        RECT 100.230 94.300 100.540 96.880 ;
        RECT 100.810 96.720 101.040 96.880 ;
        RECT 105.330 94.300 105.710 99.660 ;
        RECT 62.780 93.410 85.520 94.060 ;
        RECT 95.440 93.650 118.240 94.300 ;
        RECT 95.440 93.450 97.300 93.650 ;
        RECT 62.780 93.230 64.640 93.410 ;
        RECT 103.990 73.560 104.360 74.800 ;
        RECT 72.340 71.040 72.710 72.280 ;
        RECT 66.670 68.430 66.900 68.520 ;
        RECT 67.810 68.430 68.040 68.520 ;
        RECT 66.670 68.260 68.040 68.430 ;
        RECT 66.670 68.100 66.900 68.260 ;
        RECT 62.780 65.680 63.840 65.930 ;
        RECT 67.230 65.680 67.540 68.260 ;
        RECT 67.810 68.100 68.040 68.260 ;
        RECT 72.330 65.680 72.710 71.040 ;
        RECT 98.320 70.950 98.550 71.040 ;
        RECT 99.460 70.950 99.690 71.040 ;
        RECT 98.320 70.780 99.690 70.950 ;
        RECT 98.320 70.620 98.550 70.780 ;
        RECT 94.450 68.200 95.450 68.420 ;
        RECT 98.880 68.200 99.190 70.780 ;
        RECT 99.460 70.620 99.690 70.780 ;
        RECT 103.980 68.200 104.360 73.560 ;
        RECT 94.450 67.550 116.890 68.200 ;
        RECT 94.450 67.420 95.450 67.550 ;
        RECT 62.780 65.630 85.240 65.680 ;
        RECT 94.540 65.630 95.410 67.420 ;
        RECT 62.780 65.080 95.410 65.630 ;
        RECT 62.780 65.030 94.380 65.080 ;
        RECT 62.780 64.910 63.840 65.030 ;
        RECT 84.170 64.990 94.380 65.030 ;
        RECT 62.800 64.900 63.800 64.910 ;
        RECT 74.740 57.440 75.190 57.640 ;
        RECT 74.740 56.990 75.170 57.440 ;
        RECT 74.720 56.840 75.180 56.990 ;
        RECT 74.200 56.580 74.430 56.710 ;
        RECT 74.740 56.690 75.180 56.840 ;
        RECT 74.730 56.580 75.180 56.690 ;
        RECT 75.340 56.580 75.570 56.710 ;
        RECT 74.200 56.330 75.570 56.580 ;
        RECT 74.200 56.210 74.430 56.330 ;
        RECT 74.730 56.220 75.180 56.330 ;
        RECT 74.740 55.830 75.180 56.220 ;
        RECT 75.340 56.210 75.570 56.330 ;
        RECT 89.150 56.280 89.600 56.480 ;
        RECT 89.150 55.830 89.580 56.280 ;
        RECT 74.750 54.760 75.160 55.830 ;
        RECT 89.130 55.680 89.590 55.830 ;
        RECT 88.610 55.420 88.840 55.550 ;
        RECT 89.150 55.530 89.590 55.680 ;
        RECT 89.140 55.420 89.590 55.530 ;
        RECT 89.750 55.420 89.980 55.550 ;
        RECT 88.610 55.170 89.980 55.420 ;
        RECT 88.610 55.050 88.840 55.170 ;
        RECT 89.140 55.060 89.590 55.170 ;
        RECT 74.500 54.620 75.490 54.760 ;
        RECT 89.150 54.670 89.590 55.060 ;
        RECT 89.750 55.050 89.980 55.170 ;
        RECT 74.440 53.760 75.490 54.620 ;
        RECT 74.440 24.960 75.470 53.760 ;
        RECT 89.160 53.600 89.570 54.670 ;
        RECT 88.910 52.820 89.900 53.600 ;
        RECT 88.900 52.600 89.900 52.820 ;
        RECT 89.190 51.530 89.680 52.600 ;
        RECT 88.020 49.670 90.140 51.530 ;
        RECT 102.580 51.340 104.030 51.630 ;
        RECT 102.580 49.860 104.090 51.340 ;
        RECT 71.710 17.600 73.800 18.290 ;
        RECT 74.510 17.710 75.470 24.960 ;
        RECT 78.650 21.480 88.610 21.695 ;
        RECT 90.420 21.480 100.380 21.765 ;
        RECT 78.650 19.860 100.380 21.480 ;
        RECT 78.650 19.650 88.610 19.860 ;
        RECT 88.890 17.800 90.070 19.860 ;
        RECT 90.420 19.720 100.380 19.860 ;
        RECT 103.180 17.800 104.090 49.860 ;
        RECT 88.890 17.790 90.650 17.800 ;
        RECT 77.370 17.770 96.440 17.790 ;
        RECT 100.290 17.770 104.090 17.800 ;
        RECT 77.370 17.710 104.090 17.770 ;
        RECT 74.510 17.600 104.090 17.710 ;
        RECT 71.710 17.100 104.090 17.600 ;
        RECT 71.710 17.010 85.540 17.100 ;
        RECT 88.890 17.050 104.090 17.100 ;
        RECT 71.710 16.680 73.800 17.010 ;
        RECT 74.510 17.000 85.540 17.010 ;
        RECT 89.650 17.010 104.090 17.050 ;
        RECT 89.650 16.990 94.950 17.010 ;
        RECT 89.650 16.800 90.650 16.990 ;
        RECT 100.290 16.980 104.090 17.010 ;
      LAYER met2 ;
        RECT 101.430 204.380 101.720 204.840 ;
        RECT 101.480 203.260 101.650 204.380 ;
        RECT 101.400 202.800 101.690 203.260 ;
        RECT 101.480 202.780 101.650 202.800 ;
        RECT 77.370 199.710 79.030 201.680 ;
        RECT 101.480 201.600 101.630 202.780 ;
        RECT 101.350 201.150 101.810 201.600 ;
        RECT 62.830 93.180 64.590 94.430 ;
        RECT 95.490 93.400 97.250 94.650 ;
        RECT 62.670 64.840 63.970 66.080 ;
        RECT 88.070 51.280 90.090 51.580 ;
        RECT 102.630 51.280 103.980 51.680 ;
        RECT 88.070 50.210 103.980 51.280 ;
        RECT 88.070 49.620 90.090 50.210 ;
        RECT 102.630 49.810 103.980 50.210 ;
        RECT 71.760 16.630 73.750 18.340 ;
      LAYER met3 ;
        RECT 22.070 201.060 23.810 201.770 ;
        RECT 32.580 201.060 34.570 201.250 ;
        RECT 21.770 201.050 35.620 201.060 ;
        RECT 77.320 201.050 79.080 201.655 ;
        RECT 21.770 200.570 81.120 201.050 ;
        RECT 21.770 200.240 35.620 200.570 ;
        RECT 22.070 199.620 23.810 200.240 ;
        RECT 77.320 199.735 79.080 200.570 ;
        RECT 21.900 94.460 35.990 94.650 ;
        RECT 95.440 94.460 97.300 94.625 ;
        RECT 21.900 93.360 120.480 94.460 ;
        RECT 21.900 93.230 35.990 93.360 ;
        RECT 62.780 93.205 64.640 93.360 ;
        RECT 21.900 64.750 24.180 65.000 ;
        RECT 32.580 64.790 44.780 64.830 ;
        RECT 62.330 64.790 64.040 66.070 ;
        RECT 32.580 64.750 64.040 64.790 ;
        RECT 21.900 64.140 64.040 64.750 ;
        RECT 21.900 63.030 64.090 64.140 ;
        RECT 32.580 63.010 64.090 63.030 ;
        RECT 32.580 19.070 32.930 19.600 ;
        RECT 20.990 19.030 32.930 19.070 ;
        RECT 39.880 19.030 76.580 19.290 ;
        RECT 20.990 16.670 76.580 19.030 ;
        RECT 21.650 16.500 23.440 16.670 ;
        RECT 32.580 16.600 76.580 16.670 ;
        RECT 32.580 16.580 39.640 16.600 ;
      LAYER met4 ;
        RECT 22.050 94.655 24.050 219.660 ;
        RECT 21.945 93.225 24.050 94.655 ;
        RECT 22.050 65.005 24.050 93.225 ;
        RECT 21.945 63.025 24.135 65.005 ;
        RECT 22.050 18.715 24.050 63.025 ;
        RECT 21.695 16.495 24.050 18.715 ;
        RECT 22.050 3.900 24.050 16.495 ;
    END
    PORT
      LAYER li1 ;
        RECT 78.480 206.650 78.980 206.820 ;
        RECT 78.480 205.600 78.980 205.770 ;
      LAYER met1 ;
        RECT 78.500 206.620 78.960 206.850 ;
        RECT 80.680 205.950 81.680 206.150 ;
        RECT 84.190 205.950 85.190 206.220 ;
        RECT 78.500 205.710 78.960 205.800 ;
        RECT 80.680 205.710 85.190 205.950 ;
        RECT 78.500 205.570 85.190 205.710 ;
        RECT 78.670 205.510 85.190 205.570 ;
        RECT 80.680 205.350 85.190 205.510 ;
        RECT 80.680 205.150 81.680 205.350 ;
        RECT 84.190 205.220 85.190 205.350 ;
      LAYER met2 ;
        RECT 111.860 218.260 147.090 218.370 ;
        RECT 84.400 218.050 147.090 218.260 ;
        RECT 84.400 217.150 147.200 218.050 ;
        RECT 84.400 217.110 147.090 217.150 ;
        RECT 84.440 206.010 84.930 217.110 ;
        RECT 111.860 217.100 147.090 217.110 ;
        RECT 84.440 205.290 84.970 206.010 ;
      LAYER met3 ;
        RECT 145.830 219.000 147.410 220.220 ;
        RECT 146.090 218.025 147.140 219.000 ;
        RECT 146.040 217.175 147.250 218.025 ;
      LAYER met4 ;
        RECT 146.590 224.680 146.890 225.760 ;
        RECT 146.420 224.660 146.890 224.680 ;
        RECT 146.420 220.225 147.060 224.660 ;
        RECT 145.875 218.995 147.365 220.225 ;
    END
  END VGND
  PIN Vr
    ANTENNAGATEAREA 3.840000 ;
    PORT
      LAYER li1 ;
        RECT 73.500 102.620 75.100 102.790 ;
        RECT 73.500 100.870 75.100 101.040 ;
        RECT 73.220 74.240 74.820 74.410 ;
        RECT 73.220 72.490 74.820 72.660 ;
      LAYER met1 ;
        RECT 73.520 102.590 75.080 102.820 ;
        RECT 74.140 101.230 74.390 102.590 ;
        RECT 77.040 102.400 78.040 102.740 ;
        RECT 83.100 102.580 84.100 102.590 ;
        RECT 83.100 102.500 87.480 102.580 ;
        RECT 83.100 102.400 87.560 102.500 ;
        RECT 77.040 102.110 87.560 102.400 ;
        RECT 77.040 101.740 78.040 102.110 ;
        RECT 74.140 101.070 74.400 101.230 ;
        RECT 73.520 100.840 75.080 101.070 ;
        RECT 77.360 101.010 77.730 101.740 ;
        RECT 83.100 101.690 87.560 102.110 ;
        RECT 83.100 101.590 84.100 101.690 ;
        RECT 74.170 100.320 74.400 100.840 ;
        RECT 77.360 100.320 77.740 101.010 ;
        RECT 74.170 100.030 77.740 100.320 ;
        RECT 77.360 99.990 77.740 100.030 ;
        RECT 73.240 74.210 74.800 74.440 ;
        RECT 76.760 74.270 77.760 74.360 ;
        RECT 86.890 74.270 87.560 101.690 ;
        RECT 73.860 72.850 74.110 74.210 ;
        RECT 76.760 73.630 87.560 74.270 ;
        RECT 76.760 73.360 77.760 73.630 ;
        RECT 86.890 73.510 87.560 73.630 ;
        RECT 73.860 72.690 74.120 72.850 ;
        RECT 73.240 72.460 74.800 72.690 ;
        RECT 77.080 72.630 77.450 73.360 ;
        RECT 73.890 71.940 74.120 72.460 ;
        RECT 77.080 71.970 77.460 72.630 ;
        RECT 77.060 71.940 77.500 71.970 ;
        RECT 73.890 71.650 77.500 71.940 ;
        RECT 77.060 69.970 77.500 71.650 ;
        RECT 77.050 69.410 77.500 69.970 ;
        RECT 77.050 67.810 77.490 69.410 ;
        RECT 76.760 67.000 77.650 67.810 ;
      LAYER met2 ;
        RECT 76.810 66.950 77.600 67.860 ;
      LAYER met3 ;
        RECT 76.760 67.710 77.650 67.835 ;
        RECT 76.420 66.540 143.360 67.710 ;
        RECT 141.070 10.150 143.320 66.540 ;
        RECT 141.010 7.280 143.430 10.150 ;
      LAYER met4 ;
        RECT 141.055 8.470 143.385 10.155 ;
        RECT 141.055 7.500 152.540 8.470 ;
        RECT 141.055 7.275 143.385 7.500 ;
        RECT 151.910 1.000 152.630 7.500 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END Vr
  PIN Vin4
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER li1 ;
        RECT 58.130 171.210 58.630 171.380 ;
        RECT 58.130 168.570 58.630 168.740 ;
        RECT 58.200 166.360 58.700 166.530 ;
        RECT 58.200 164.810 58.700 164.980 ;
      LAYER met1 ;
        RECT 58.150 171.180 58.610 171.410 ;
        RECT 58.150 168.540 58.610 168.770 ;
        RECT 54.050 167.810 55.050 168.040 ;
        RECT 55.330 167.810 56.330 168.080 ;
        RECT 58.300 167.810 58.440 168.540 ;
        RECT 54.050 167.530 58.460 167.810 ;
        RECT 54.050 167.040 55.050 167.530 ;
        RECT 55.330 167.080 56.330 167.530 ;
        RECT 58.300 166.560 58.440 167.530 ;
        RECT 58.220 166.330 58.680 166.560 ;
        RECT 58.220 164.780 58.680 165.010 ;
      LAYER met2 ;
        RECT 54.160 167.990 54.820 168.040 ;
        RECT 54.120 167.090 54.830 167.990 ;
        RECT 55.400 167.200 56.100 168.030 ;
      LAYER met3 ;
        RECT 119.810 212.140 121.430 212.180 ;
        RECT 119.730 210.210 121.430 212.140 ;
        RECT 119.810 195.710 121.430 210.210 ;
        RECT 56.530 195.640 121.570 195.710 ;
        RECT 54.020 194.680 121.570 195.640 ;
        RECT 54.020 194.460 60.450 194.680 ;
        RECT 54.020 167.965 54.840 194.460 ;
        RECT 54.020 167.910 54.880 167.965 ;
        RECT 55.350 167.910 56.150 168.005 ;
        RECT 54.020 167.225 56.150 167.910 ;
        RECT 54.020 167.160 56.050 167.225 ;
        RECT 54.020 167.115 54.880 167.160 ;
        RECT 54.020 166.990 54.840 167.115 ;
      LAYER met4 ;
        RECT 130.030 224.670 130.330 225.760 ;
        RECT 130.020 223.590 130.330 224.670 ;
        RECT 119.840 222.800 130.330 223.590 ;
        RECT 119.840 222.780 129.630 222.800 ;
        RECT 119.840 212.145 121.080 222.780 ;
        RECT 119.775 210.205 121.355 212.145 ;
    END
  END Vin4
  PIN Vin3
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER li1 ;
        RECT 76.640 170.600 77.140 170.770 ;
        RECT 76.640 167.960 77.140 168.130 ;
        RECT 76.710 165.750 77.210 165.920 ;
        RECT 76.710 164.200 77.210 164.370 ;
      LAYER met1 ;
        RECT 76.660 170.570 77.120 170.800 ;
        RECT 76.660 167.930 77.120 168.160 ;
        RECT 69.690 167.260 70.690 167.530 ;
        RECT 72.560 167.260 73.560 167.430 ;
        RECT 69.690 167.200 73.560 167.260 ;
        RECT 76.810 167.200 76.950 167.930 ;
        RECT 69.690 166.920 76.970 167.200 ;
        RECT 69.690 166.800 73.560 166.920 ;
        RECT 69.690 166.530 70.690 166.800 ;
        RECT 72.560 166.430 73.560 166.800 ;
        RECT 76.810 165.950 76.950 166.920 ;
        RECT 76.730 165.720 77.190 165.950 ;
        RECT 76.730 164.170 77.190 164.400 ;
      LAYER met2 ;
        RECT 69.780 166.550 70.550 167.460 ;
      LAYER met3 ;
        RECT 123.600 210.060 125.270 211.990 ;
        RECT 69.960 193.740 70.840 193.890 ;
        RECT 69.820 193.670 86.370 193.740 ;
        RECT 124.050 193.670 124.870 210.060 ;
        RECT 69.820 192.710 125.050 193.670 ;
        RECT 69.960 167.435 70.840 192.710 ;
        RECT 79.710 192.570 125.050 192.710 ;
        RECT 124.050 192.480 124.870 192.570 ;
        RECT 69.730 166.575 70.840 167.435 ;
        RECT 69.960 166.490 70.840 166.575 ;
      LAYER met4 ;
        RECT 132.790 224.670 133.090 225.760 ;
        RECT 132.770 224.390 133.090 224.670 ;
        RECT 132.760 223.690 133.070 224.390 ;
        RECT 124.010 221.580 124.750 221.610 ;
        RECT 132.750 221.580 133.080 223.690 ;
        RECT 124.010 221.560 133.090 221.580 ;
        RECT 124.010 220.780 133.150 221.560 ;
        RECT 124.010 220.770 133.090 220.780 ;
        RECT 124.010 211.995 124.750 220.770 ;
        RECT 123.645 210.055 125.225 211.995 ;
    END
    PORT
      LAYER li1 ;
        RECT 82.410 40.255 82.580 40.795 ;
        RECT 78.630 33.650 88.630 33.820 ;
        RECT 78.710 31.835 88.550 33.650 ;
      LAYER met1 ;
        RECT 82.380 40.610 82.610 40.775 ;
        RECT 82.380 40.275 82.810 40.610 ;
        RECT 77.330 37.820 78.330 38.200 ;
        RECT 80.180 37.880 81.180 38.190 ;
        RECT 82.500 37.880 82.810 40.275 ;
        RECT 80.180 37.820 82.810 37.880 ;
        RECT 77.330 37.350 82.810 37.820 ;
        RECT 77.330 37.200 78.330 37.350 ;
        RECT 80.180 37.310 82.810 37.350 ;
        RECT 80.180 37.190 81.180 37.310 ;
        RECT 82.010 33.850 82.320 33.890 ;
        RECT 82.500 33.850 82.810 37.310 ;
        RECT 78.650 31.805 88.610 33.850 ;
      LAYER met2 ;
        RECT 62.840 38.150 64.440 38.220 ;
        RECT 62.840 38.040 78.040 38.150 ;
        RECT 62.840 37.390 78.100 38.040 ;
        RECT 62.840 37.160 78.040 37.390 ;
        RECT 62.840 12.630 64.440 37.160 ;
        RECT 125.950 12.630 127.880 12.680 ;
        RECT 62.710 11.160 127.880 12.630 ;
        RECT 62.710 11.040 127.430 11.160 ;
      LAYER met3 ;
        RECT 125.900 12.630 127.930 12.655 ;
        RECT 132.080 12.630 133.770 12.740 ;
        RECT 125.900 11.210 133.770 12.630 ;
        RECT 125.900 11.185 127.930 11.210 ;
        RECT 132.080 11.040 133.770 11.210 ;
      LAYER met4 ;
        RECT 132.125 11.035 133.725 12.745 ;
        RECT 132.360 8.600 133.320 11.035 ;
        RECT 132.560 1.000 133.280 8.600 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END Vin3
  PIN Vin2
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER li1 ;
        RECT 99.110 171.130 99.610 171.300 ;
        RECT 99.110 168.490 99.610 168.660 ;
        RECT 99.180 166.280 99.680 166.450 ;
        RECT 99.180 164.730 99.680 164.900 ;
      LAYER met1 ;
        RECT 99.130 171.100 99.590 171.330 ;
        RECT 99.130 168.460 99.590 168.690 ;
        RECT 92.810 167.850 93.810 167.960 ;
        RECT 92.810 167.640 93.850 167.850 ;
        RECT 95.030 167.730 96.030 167.960 ;
        RECT 99.280 167.730 99.420 168.460 ;
        RECT 95.030 167.640 99.440 167.730 ;
        RECT 92.810 167.450 99.440 167.640 ;
        RECT 92.810 167.190 96.030 167.450 ;
        RECT 92.810 167.180 93.850 167.190 ;
        RECT 92.810 166.960 93.810 167.180 ;
        RECT 95.030 166.960 96.030 167.190 ;
        RECT 99.280 166.480 99.420 167.450 ;
        RECT 99.200 166.250 99.660 166.480 ;
        RECT 99.200 164.700 99.660 164.930 ;
      LAYER met2 ;
        RECT 93.050 167.130 93.800 167.900 ;
      LAYER met3 ;
        RECT 126.890 209.710 128.560 211.640 ;
        RECT 93.110 192.100 93.910 192.180 ;
        RECT 93.110 191.880 95.450 192.100 ;
        RECT 127.390 191.920 128.010 209.710 ;
        RECT 108.840 191.880 128.010 191.920 ;
        RECT 93.110 191.300 128.010 191.880 ;
        RECT 93.110 167.875 93.910 191.300 ;
        RECT 108.840 191.250 128.010 191.300 ;
        RECT 93.000 167.380 93.910 167.875 ;
        RECT 93.000 167.155 93.850 167.380 ;
      LAYER met4 ;
        RECT 135.550 224.300 135.850 225.760 ;
        RECT 135.490 220.180 135.880 224.300 ;
        RECT 129.470 220.170 135.900 220.180 ;
        RECT 127.260 219.660 135.900 220.170 ;
        RECT 127.260 219.530 130.440 219.660 ;
        RECT 127.330 211.645 128.070 219.530 ;
        RECT 126.935 209.705 128.515 211.645 ;
    END
    PORT
      LAYER li1 ;
        RECT 83.550 40.255 83.720 40.795 ;
        RECT 90.400 33.720 100.400 33.890 ;
        RECT 90.480 31.905 100.320 33.720 ;
      LAYER met1 ;
        RECT 83.520 40.730 83.750 40.775 ;
        RECT 83.440 40.275 83.750 40.730 ;
        RECT 83.440 38.010 83.640 40.275 ;
        RECT 84.680 38.010 85.680 38.320 ;
        RECT 83.440 37.920 85.680 38.010 ;
        RECT 87.650 37.920 88.650 38.290 ;
        RECT 83.440 37.650 88.650 37.920 ;
        RECT 83.440 37.440 85.680 37.650 ;
        RECT 83.440 36.010 83.640 37.440 ;
        RECT 84.680 37.320 85.680 37.440 ;
        RECT 87.650 37.290 88.650 37.650 ;
        RECT 86.690 36.010 93.890 36.050 ;
        RECT 95.370 36.010 95.760 36.040 ;
        RECT 83.440 35.700 95.760 36.010 ;
        RECT 83.950 35.680 95.760 35.700 ;
        RECT 86.690 35.650 93.890 35.680 ;
        RECT 95.370 33.920 95.760 35.680 ;
        RECT 90.420 31.875 100.380 33.920 ;
      LAYER met2 ;
        RECT 112.640 38.190 113.470 38.210 ;
        RECT 109.940 38.150 114.250 38.190 ;
        RECT 87.710 37.600 114.250 38.150 ;
        RECT 87.780 37.440 88.360 37.600 ;
        RECT 109.640 37.520 114.250 37.600 ;
        RECT 109.640 37.490 110.780 37.520 ;
        RECT 112.640 37.500 113.470 37.520 ;
      LAYER met3 ;
        RECT 112.590 38.170 113.520 38.185 ;
        RECT 112.580 36.540 113.560 38.170 ;
        RECT 112.560 10.810 113.610 36.540 ;
        RECT 112.130 8.600 114.550 10.810 ;
      LAYER met4 ;
        RECT 112.175 8.595 114.505 10.815 ;
        RECT 113.280 1.000 114.000 8.595 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END Vin2
  PIN Vin1
    ANTENNAGATEAREA 1.500000 ;
    PORT
      LAYER li1 ;
        RECT 114.690 158.150 115.190 158.320 ;
        RECT 114.690 155.510 115.190 155.680 ;
        RECT 114.760 153.300 115.260 153.470 ;
        RECT 114.760 151.750 115.260 151.920 ;
      LAYER met1 ;
        RECT 114.710 158.120 115.170 158.350 ;
        RECT 114.710 155.480 115.170 155.710 ;
        RECT 108.450 154.870 109.450 154.960 ;
        RECT 110.610 154.870 111.610 154.980 ;
        RECT 108.450 154.750 111.620 154.870 ;
        RECT 114.860 154.750 115.000 155.480 ;
        RECT 108.450 154.470 115.020 154.750 ;
        RECT 108.450 154.160 111.620 154.470 ;
        RECT 108.450 153.960 109.450 154.160 ;
        RECT 110.610 153.980 111.610 154.160 ;
        RECT 114.860 153.500 115.000 154.470 ;
        RECT 114.780 153.270 115.240 153.500 ;
        RECT 114.780 151.720 115.240 151.950 ;
      LAYER met2 ;
        RECT 108.630 153.970 109.390 154.890 ;
      LAYER met3 ;
        RECT 128.960 209.780 130.630 211.710 ;
        RECT 129.190 201.920 130.300 209.780 ;
        RECT 108.790 190.480 109.510 190.560 ;
        RECT 128.900 190.480 130.570 201.920 ;
        RECT 108.720 189.110 130.710 190.480 ;
        RECT 108.790 154.865 109.510 189.110 ;
        RECT 108.580 154.020 109.510 154.865 ;
        RECT 108.580 153.995 109.440 154.020 ;
      LAYER met4 ;
        RECT 138.310 223.650 138.610 225.760 ;
        RECT 138.280 222.380 138.610 223.650 ;
        RECT 130.350 218.940 137.740 218.960 ;
        RECT 138.170 218.940 138.670 222.380 ;
        RECT 130.350 218.860 138.670 218.940 ;
        RECT 129.410 218.310 138.670 218.860 ;
        RECT 129.410 218.300 136.610 218.310 ;
        RECT 129.410 211.715 130.040 218.300 ;
        RECT 129.005 209.775 130.585 211.715 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END Vin1
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.380 224.660 49.680 225.660 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 57.220 164.120 59.680 167.220 ;
        RECT 75.730 163.510 78.190 166.610 ;
        RECT 98.200 164.040 100.660 167.140 ;
        RECT 45.850 154.650 49.290 161.180 ;
        RECT 66.190 158.240 68.650 161.340 ;
        RECT 88.720 159.020 91.180 162.120 ;
        RECT 109.660 159.510 112.120 162.610 ;
        RECT 127.090 159.180 129.550 162.280 ;
        RECT 96.730 146.820 99.390 154.430 ;
        RECT 100.820 146.700 103.480 154.310 ;
        RECT 113.780 151.060 116.240 154.160 ;
        RECT 77.800 18.770 89.460 34.730 ;
        RECT 89.570 18.840 101.230 34.800 ;
      LAYER li1 ;
        RECT 94.890 212.400 96.490 212.570 ;
        RECT 96.780 212.400 98.380 212.570 ;
        RECT 99.810 212.400 101.410 212.570 ;
        RECT 101.700 212.400 103.300 212.570 ;
        RECT 94.660 211.725 94.830 212.185 ;
        RECT 98.440 211.725 98.610 212.185 ;
        RECT 99.580 211.725 99.750 212.185 ;
        RECT 101.470 211.725 101.640 212.185 ;
        RECT 103.360 211.725 103.530 212.185 ;
        RECT 94.890 211.340 96.490 211.510 ;
        RECT 96.780 211.340 98.380 211.510 ;
        RECT 99.810 211.340 101.410 211.510 ;
        RECT 101.700 211.340 103.300 211.510 ;
        RECT 94.890 210.800 96.490 210.970 ;
        RECT 96.780 210.800 98.380 210.970 ;
        RECT 99.810 210.800 101.410 210.970 ;
        RECT 101.700 210.800 103.300 210.970 ;
        RECT 94.660 210.125 94.830 210.585 ;
        RECT 98.440 210.125 98.610 210.585 ;
        RECT 99.580 210.125 99.750 210.585 ;
        RECT 101.470 210.125 101.640 210.585 ;
        RECT 103.360 210.125 103.530 210.585 ;
        RECT 78.460 209.790 78.960 209.960 ;
        RECT 94.890 209.740 96.490 209.910 ;
        RECT 96.780 209.740 98.380 209.910 ;
        RECT 99.810 209.740 101.410 209.910 ;
        RECT 101.700 209.740 103.300 209.910 ;
        RECT 73.990 209.070 74.990 209.240 ;
        RECT 79.020 209.035 79.190 209.575 ;
        RECT 73.760 207.815 73.930 208.855 ;
        RECT 78.460 208.650 78.960 208.820 ;
        RECT 94.890 208.720 96.490 208.890 ;
        RECT 96.780 208.720 98.380 208.890 ;
        RECT 99.810 208.720 101.410 208.890 ;
        RECT 101.700 208.720 103.300 208.890 ;
        RECT 94.660 208.045 94.830 208.505 ;
        RECT 96.550 208.045 96.720 208.505 ;
        RECT 98.440 208.045 98.610 208.505 ;
        RECT 99.580 208.045 99.750 208.505 ;
        RECT 101.470 208.045 101.640 208.505 ;
        RECT 103.360 208.045 103.530 208.505 ;
        RECT 94.890 207.660 96.490 207.830 ;
        RECT 96.780 207.660 98.380 207.830 ;
        RECT 99.810 207.660 101.410 207.830 ;
        RECT 101.700 207.660 103.300 207.830 ;
        RECT 73.990 207.430 74.990 207.600 ;
        RECT 94.890 207.120 96.490 207.290 ;
        RECT 96.780 207.120 98.380 207.290 ;
        RECT 99.810 207.120 101.410 207.290 ;
        RECT 101.700 207.120 103.300 207.290 ;
        RECT 73.990 206.890 74.990 207.060 ;
        RECT 73.760 205.635 73.930 206.675 ;
        RECT 79.040 205.940 79.210 206.480 ;
        RECT 94.660 206.445 94.830 206.905 ;
        RECT 96.550 206.445 96.720 206.905 ;
        RECT 98.440 206.445 98.610 206.905 ;
        RECT 99.580 206.445 99.750 206.905 ;
        RECT 101.470 206.445 101.640 206.905 ;
        RECT 103.360 206.445 103.530 206.905 ;
        RECT 94.890 206.060 96.490 206.230 ;
        RECT 96.780 206.060 98.380 206.230 ;
        RECT 99.810 206.060 101.410 206.230 ;
        RECT 101.700 206.060 103.300 206.230 ;
        RECT 73.990 205.250 74.990 205.420 ;
        RECT 94.890 205.040 96.490 205.210 ;
        RECT 96.780 205.040 98.380 205.210 ;
        RECT 94.660 204.365 94.830 204.825 ;
        RECT 96.550 204.365 96.720 204.825 ;
        RECT 98.440 204.365 98.610 204.825 ;
        RECT 99.580 204.365 99.750 204.825 ;
        RECT 103.360 204.365 103.530 204.825 ;
        RECT 94.890 203.980 96.490 204.150 ;
        RECT 96.780 203.980 98.380 204.150 ;
        RECT 94.890 203.440 96.490 203.610 ;
        RECT 96.780 203.440 98.380 203.610 ;
        RECT 94.660 202.765 94.830 203.225 ;
        RECT 96.550 202.765 96.720 203.225 ;
        RECT 98.440 202.765 98.610 203.225 ;
        RECT 99.580 202.765 99.750 203.225 ;
        RECT 103.360 202.765 103.530 203.225 ;
        RECT 94.890 202.380 96.490 202.550 ;
        RECT 96.780 202.380 98.380 202.550 ;
        RECT 67.415 183.080 67.745 183.250 ;
        RECT 68.005 183.080 68.335 183.250 ;
        RECT 69.735 183.080 70.065 183.250 ;
        RECT 70.325 183.080 70.655 183.250 ;
        RECT 46.755 180.600 47.085 180.770 ;
        RECT 47.345 180.600 47.675 180.770 ;
        RECT 47.935 180.600 48.265 180.770 ;
        RECT 46.540 179.925 46.710 180.385 ;
        RECT 47.720 179.925 47.890 180.385 ;
        RECT 67.790 180.325 67.960 182.865 ;
        RECT 70.110 180.325 70.280 182.865 ;
        RECT 109.615 182.730 109.945 182.900 ;
        RECT 110.205 182.730 110.535 182.900 ;
        RECT 111.935 182.730 112.265 182.900 ;
        RECT 112.525 182.730 112.855 182.900 ;
        RECT 89.835 182.400 90.165 182.570 ;
        RECT 90.425 182.400 90.755 182.570 ;
        RECT 92.155 182.400 92.485 182.570 ;
        RECT 92.745 182.400 93.075 182.570 ;
        RECT 67.415 179.940 67.745 180.110 ;
        RECT 68.005 179.940 68.335 180.110 ;
        RECT 69.735 179.940 70.065 180.110 ;
        RECT 70.325 179.940 70.655 180.110 ;
        RECT 46.755 179.540 47.085 179.710 ;
        RECT 47.345 179.540 47.675 179.710 ;
        RECT 47.935 179.540 48.265 179.710 ;
        RECT 89.620 179.645 89.790 182.185 ;
        RECT 90.210 179.645 90.380 182.185 ;
        RECT 90.800 179.645 90.970 182.185 ;
        RECT 91.940 179.645 92.110 182.185 ;
        RECT 92.530 179.645 92.700 182.185 ;
        RECT 93.120 179.645 93.290 182.185 ;
        RECT 109.400 179.975 109.570 182.515 ;
        RECT 109.990 179.975 110.160 182.515 ;
        RECT 110.580 179.975 110.750 182.515 ;
        RECT 111.720 179.975 111.890 182.515 ;
        RECT 112.310 179.975 112.480 182.515 ;
        RECT 112.900 179.975 113.070 182.515 ;
        RECT 128.645 181.730 128.975 181.900 ;
        RECT 129.235 181.730 129.565 181.900 ;
        RECT 109.615 179.590 109.945 179.760 ;
        RECT 110.205 179.590 110.535 179.760 ;
        RECT 111.935 179.590 112.265 179.760 ;
        RECT 112.525 179.590 112.855 179.760 ;
        RECT 89.835 179.260 90.165 179.430 ;
        RECT 90.425 179.260 90.755 179.430 ;
        RECT 92.155 179.260 92.485 179.430 ;
        RECT 92.745 179.260 93.075 179.430 ;
        RECT 46.755 179.000 47.085 179.170 ;
        RECT 47.345 179.000 47.675 179.170 ;
        RECT 47.935 179.000 48.265 179.170 ;
        RECT 67.415 178.920 67.745 179.090 ;
        RECT 68.005 178.920 68.335 179.090 ;
        RECT 69.735 178.920 70.065 179.090 ;
        RECT 70.325 178.920 70.655 179.090 ;
        RECT 128.430 178.975 128.600 181.515 ;
        RECT 129.020 178.975 129.190 181.515 ;
        RECT 129.610 178.975 129.780 181.515 ;
        RECT 46.540 178.325 46.710 178.785 ;
        RECT 47.720 178.325 47.890 178.785 ;
        RECT 46.755 177.940 47.085 178.110 ;
        RECT 47.345 177.940 47.675 178.110 ;
        RECT 47.935 177.940 48.265 178.110 ;
        RECT 46.755 177.400 47.085 177.570 ;
        RECT 47.345 177.400 47.675 177.570 ;
        RECT 47.935 177.400 48.265 177.570 ;
        RECT 46.540 176.725 46.710 177.185 ;
        RECT 47.720 176.725 47.890 177.185 ;
        RECT 46.755 176.340 47.085 176.510 ;
        RECT 47.345 176.340 47.675 176.510 ;
        RECT 47.935 176.340 48.265 176.510 ;
        RECT 67.200 176.165 67.370 178.705 ;
        RECT 67.790 176.165 67.960 178.705 ;
        RECT 68.380 176.165 68.550 178.705 ;
        RECT 69.520 176.165 69.690 178.705 ;
        RECT 70.110 176.165 70.280 178.705 ;
        RECT 70.700 176.165 70.870 178.705 ;
        RECT 109.615 178.570 109.945 178.740 ;
        RECT 110.205 178.570 110.535 178.740 ;
        RECT 111.935 178.570 112.265 178.740 ;
        RECT 112.525 178.570 112.855 178.740 ;
        RECT 128.645 178.590 128.975 178.760 ;
        RECT 129.235 178.590 129.565 178.760 ;
        RECT 89.835 178.240 90.165 178.410 ;
        RECT 90.425 178.240 90.755 178.410 ;
        RECT 92.155 178.240 92.485 178.410 ;
        RECT 92.745 178.240 93.075 178.410 ;
        RECT 140.365 178.370 140.695 178.540 ;
        RECT 140.955 178.370 141.285 178.540 ;
        RECT 46.755 175.800 47.085 175.970 ;
        RECT 47.345 175.800 47.675 175.970 ;
        RECT 47.935 175.800 48.265 175.970 ;
        RECT 67.415 175.780 67.745 175.950 ;
        RECT 68.005 175.780 68.335 175.950 ;
        RECT 69.735 175.780 70.065 175.950 ;
        RECT 70.325 175.780 70.655 175.950 ;
        RECT 46.540 175.125 46.710 175.585 ;
        RECT 47.720 175.125 47.890 175.585 ;
        RECT 89.620 175.485 89.790 178.025 ;
        RECT 90.210 175.485 90.380 178.025 ;
        RECT 90.800 175.485 90.970 178.025 ;
        RECT 91.940 175.485 92.110 178.025 ;
        RECT 92.530 175.485 92.700 178.025 ;
        RECT 93.120 175.485 93.290 178.025 ;
        RECT 109.400 175.815 109.570 178.355 ;
        RECT 109.990 175.815 110.160 178.355 ;
        RECT 110.580 175.815 110.750 178.355 ;
        RECT 111.720 175.815 111.890 178.355 ;
        RECT 112.310 175.815 112.480 178.355 ;
        RECT 112.900 175.815 113.070 178.355 ;
        RECT 127.305 175.750 127.635 175.920 ;
        RECT 127.895 175.750 128.225 175.920 ;
        RECT 129.625 175.750 129.955 175.920 ;
        RECT 130.215 175.750 130.545 175.920 ;
        RECT 140.150 175.615 140.320 178.155 ;
        RECT 140.740 175.615 140.910 178.155 ;
        RECT 141.330 175.615 141.500 178.155 ;
        RECT 109.615 175.430 109.945 175.600 ;
        RECT 110.205 175.430 110.535 175.600 ;
        RECT 111.935 175.430 112.265 175.600 ;
        RECT 112.525 175.430 112.855 175.600 ;
        RECT 89.835 175.100 90.165 175.270 ;
        RECT 90.425 175.100 90.755 175.270 ;
        RECT 92.155 175.100 92.485 175.270 ;
        RECT 92.745 175.100 93.075 175.270 ;
        RECT 46.755 174.740 47.085 174.910 ;
        RECT 47.345 174.740 47.675 174.910 ;
        RECT 47.935 174.740 48.265 174.910 ;
        RECT 46.755 174.200 47.085 174.370 ;
        RECT 47.345 174.200 47.675 174.370 ;
        RECT 47.935 174.200 48.265 174.370 ;
        RECT 46.540 173.525 46.710 173.985 ;
        RECT 47.720 173.525 47.890 173.985 ;
        RECT 46.755 173.140 47.085 173.310 ;
        RECT 47.345 173.140 47.675 173.310 ;
        RECT 47.935 173.140 48.265 173.310 ;
        RECT 127.090 172.995 127.260 175.535 ;
        RECT 127.680 172.995 127.850 175.535 ;
        RECT 128.270 172.995 128.440 175.535 ;
        RECT 129.410 172.995 129.580 175.535 ;
        RECT 130.000 172.995 130.170 175.535 ;
        RECT 130.590 172.995 130.760 175.535 ;
        RECT 140.365 175.230 140.695 175.400 ;
        RECT 140.955 175.230 141.285 175.400 ;
        RECT 46.755 172.600 47.085 172.770 ;
        RECT 47.345 172.600 47.675 172.770 ;
        RECT 47.935 172.600 48.265 172.770 ;
        RECT 127.305 172.610 127.635 172.780 ;
        RECT 127.895 172.610 128.225 172.780 ;
        RECT 129.625 172.610 129.955 172.780 ;
        RECT 130.215 172.610 130.545 172.780 ;
        RECT 46.540 171.925 46.710 172.385 ;
        RECT 47.720 171.925 47.890 172.385 ;
        RECT 46.755 171.540 47.085 171.710 ;
        RECT 47.345 171.540 47.675 171.710 ;
        RECT 47.935 171.540 48.265 171.710 ;
        RECT 46.755 171.000 47.085 171.170 ;
        RECT 47.345 171.000 47.675 171.170 ;
        RECT 47.935 171.000 48.265 171.170 ;
        RECT 46.540 170.325 46.710 170.785 ;
        RECT 47.720 170.325 47.890 170.785 ;
        RECT 46.755 169.940 47.085 170.110 ;
        RECT 47.345 169.940 47.675 170.110 ;
        RECT 47.935 169.940 48.265 170.110 ;
        RECT 46.755 169.400 47.085 169.570 ;
        RECT 47.345 169.400 47.675 169.570 ;
        RECT 47.935 169.400 48.265 169.570 ;
        RECT 46.540 168.725 46.710 169.185 ;
        RECT 47.720 168.725 47.890 169.185 ;
        RECT 58.690 168.955 58.860 170.995 ;
        RECT 46.755 168.340 47.085 168.510 ;
        RECT 47.345 168.340 47.675 168.510 ;
        RECT 47.935 168.340 48.265 168.510 ;
        RECT 77.200 168.345 77.370 170.385 ;
        RECT 99.670 168.875 99.840 170.915 ;
        RECT 46.755 167.800 47.085 167.970 ;
        RECT 47.345 167.800 47.675 167.970 ;
        RECT 47.935 167.800 48.265 167.970 ;
        RECT 46.540 167.125 46.710 167.585 ;
        RECT 47.720 167.125 47.890 167.585 ;
        RECT 46.755 166.740 47.085 166.910 ;
        RECT 47.345 166.740 47.675 166.910 ;
        RECT 47.935 166.740 48.265 166.910 ;
        RECT 57.400 166.870 59.500 167.040 ;
        RECT 46.755 166.200 47.085 166.370 ;
        RECT 47.345 166.200 47.675 166.370 ;
        RECT 47.935 166.200 48.265 166.370 ;
        RECT 46.540 165.525 46.710 165.985 ;
        RECT 47.720 165.525 47.890 165.985 ;
        RECT 57.400 165.610 57.570 166.870 ;
        RECT 57.400 165.370 57.720 165.610 ;
        RECT 46.755 165.140 47.085 165.310 ;
        RECT 47.345 165.140 47.675 165.310 ;
        RECT 47.935 165.140 48.265 165.310 ;
        RECT 57.400 164.470 57.570 165.370 ;
        RECT 57.970 165.150 58.140 166.190 ;
        RECT 58.760 165.150 58.930 166.190 ;
        RECT 59.330 164.470 59.500 166.870 ;
        RECT 98.380 166.790 100.480 166.960 ;
        RECT 75.910 166.260 78.010 166.430 ;
        RECT 67.100 165.330 67.600 165.500 ;
        RECT 57.400 164.300 59.500 164.470 ;
        RECT 67.660 163.075 67.830 165.115 ;
        RECT 75.910 165.000 76.080 166.260 ;
        RECT 75.910 164.760 76.230 165.000 ;
        RECT 75.910 163.860 76.080 164.760 ;
        RECT 76.480 164.540 76.650 165.580 ;
        RECT 77.270 164.540 77.440 165.580 ;
        RECT 77.840 163.860 78.010 166.260 ;
        RECT 89.630 166.110 90.130 166.280 ;
        RECT 75.910 163.690 78.010 163.860 ;
        RECT 90.190 163.855 90.360 165.895 ;
        RECT 98.380 165.530 98.550 166.790 ;
        RECT 98.380 165.290 98.700 165.530 ;
        RECT 98.380 164.390 98.550 165.290 ;
        RECT 98.950 165.070 99.120 166.110 ;
        RECT 99.740 165.070 99.910 166.110 ;
        RECT 100.310 164.390 100.480 166.790 ;
        RECT 110.570 166.600 111.070 166.770 ;
        RECT 98.380 164.220 100.480 164.390 ;
        RECT 111.130 164.345 111.300 166.385 ;
        RECT 128.000 166.270 128.500 166.440 ;
        RECT 110.570 163.960 111.070 164.130 ;
        RECT 128.560 164.015 128.730 166.055 ;
        RECT 140.815 165.630 141.145 165.800 ;
        RECT 141.405 165.630 141.735 165.800 ;
        RECT 89.630 163.470 90.130 163.640 ;
        RECT 128.000 163.630 128.500 163.800 ;
        RECT 140.600 162.875 140.770 165.415 ;
        RECT 141.190 162.875 141.360 165.415 ;
        RECT 141.780 162.875 141.950 165.415 ;
        RECT 67.100 162.690 67.600 162.860 ;
        RECT 140.815 162.490 141.145 162.660 ;
        RECT 141.405 162.490 141.735 162.660 ;
        RECT 109.840 162.260 111.940 162.430 ;
        RECT 88.900 161.770 91.000 161.940 ;
        RECT 46.030 160.830 49.110 161.000 ;
        RECT 46.030 155.000 46.200 160.830 ;
        RECT 46.600 158.440 46.770 160.150 ;
        RECT 47.190 158.440 47.360 160.150 ;
        RECT 47.780 158.440 47.950 160.150 ;
        RECT 48.370 158.440 48.540 160.150 ;
        RECT 46.600 155.680 46.770 157.390 ;
        RECT 47.190 155.680 47.360 157.390 ;
        RECT 47.780 155.680 47.950 157.390 ;
        RECT 48.370 155.680 48.540 157.390 ;
        RECT 48.560 155.000 48.730 155.060 ;
        RECT 48.940 155.000 49.110 160.830 ;
        RECT 66.370 160.990 68.470 161.160 ;
        RECT 66.370 159.730 66.540 160.990 ;
        RECT 67.170 160.480 67.670 160.650 ;
        RECT 66.370 159.490 66.690 159.730 ;
        RECT 66.370 158.590 66.540 159.490 ;
        RECT 66.940 159.270 67.110 160.310 ;
        RECT 67.730 159.270 67.900 160.310 ;
        RECT 67.170 158.930 67.670 159.100 ;
        RECT 68.300 158.590 68.470 160.990 ;
        RECT 88.900 160.510 89.070 161.770 ;
        RECT 89.700 161.260 90.200 161.430 ;
        RECT 88.900 160.270 89.220 160.510 ;
        RECT 88.900 159.370 89.070 160.270 ;
        RECT 89.470 160.050 89.640 161.090 ;
        RECT 90.260 160.050 90.430 161.090 ;
        RECT 89.700 159.710 90.200 159.880 ;
        RECT 90.830 159.370 91.000 161.770 ;
        RECT 109.840 161.000 110.010 162.260 ;
        RECT 110.640 161.750 111.140 161.920 ;
        RECT 109.840 160.760 110.160 161.000 ;
        RECT 109.840 159.860 110.010 160.760 ;
        RECT 110.410 160.540 110.580 161.580 ;
        RECT 111.200 160.540 111.370 161.580 ;
        RECT 110.640 160.200 111.140 160.370 ;
        RECT 111.770 159.860 111.940 162.260 ;
        RECT 109.840 159.690 111.940 159.860 ;
        RECT 127.270 161.930 129.370 162.100 ;
        RECT 127.270 160.670 127.440 161.930 ;
        RECT 128.070 161.420 128.570 161.590 ;
        RECT 127.270 160.430 127.590 160.670 ;
        RECT 88.900 159.200 91.000 159.370 ;
        RECT 127.270 159.530 127.440 160.430 ;
        RECT 127.840 160.210 128.010 161.250 ;
        RECT 128.630 160.210 128.800 161.250 ;
        RECT 128.070 159.870 128.570 160.040 ;
        RECT 129.200 159.530 129.370 161.930 ;
        RECT 127.270 159.360 129.370 159.530 ;
        RECT 66.370 158.420 68.470 158.590 ;
        RECT 115.250 155.895 115.420 157.935 ;
        RECT 46.030 154.830 49.110 155.000 ;
        RECT 96.910 154.080 99.210 154.250 ;
        RECT 96.910 147.170 97.080 154.080 ;
        RECT 97.560 153.350 98.560 153.520 ;
        RECT 97.640 151.535 98.480 153.350 ;
        RECT 97.640 147.900 98.480 149.715 ;
        RECT 99.040 148.270 99.210 154.080 ;
        RECT 101.000 153.960 103.300 154.130 ;
        RECT 99.040 147.930 99.260 148.270 ;
        RECT 97.560 147.730 98.560 147.900 ;
        RECT 99.040 147.170 99.210 147.930 ;
        RECT 96.910 147.000 99.210 147.170 ;
        RECT 101.000 147.050 101.170 153.960 ;
        RECT 101.650 153.230 102.650 153.400 ;
        RECT 101.730 151.415 102.570 153.230 ;
        RECT 101.730 147.780 102.570 149.595 ;
        RECT 103.130 148.250 103.300 153.960 ;
        RECT 113.960 153.810 116.060 153.980 ;
        RECT 113.960 152.550 114.130 153.810 ;
        RECT 113.960 152.310 114.280 152.550 ;
        RECT 113.960 151.410 114.130 152.310 ;
        RECT 114.530 152.090 114.700 153.130 ;
        RECT 115.320 152.090 115.490 153.130 ;
        RECT 115.890 151.410 116.060 153.810 ;
        RECT 113.960 151.240 116.060 151.410 ;
        RECT 103.110 147.910 103.330 148.250 ;
        RECT 101.650 147.610 102.650 147.780 ;
        RECT 103.130 147.050 103.300 147.910 ;
        RECT 101.000 146.880 103.300 147.050 ;
        RECT 111.280 112.060 112.880 112.230 ;
        RECT 114.310 112.060 115.910 112.230 ;
        RECT 78.560 111.820 80.160 111.990 ;
        RECT 81.590 111.820 83.190 111.990 ;
        RECT 97.230 111.860 98.830 112.030 ;
        RECT 100.260 111.860 101.860 112.030 ;
        RECT 64.510 111.620 66.110 111.790 ;
        RECT 67.540 111.620 69.140 111.790 ;
        RECT 64.280 110.865 64.450 111.405 ;
        RECT 69.200 110.865 69.370 111.405 ;
        RECT 78.330 111.065 78.500 111.605 ;
        RECT 83.250 111.065 83.420 111.605 ;
        RECT 97.000 111.105 97.170 111.645 ;
        RECT 101.920 111.105 102.090 111.645 ;
        RECT 111.050 111.305 111.220 111.845 ;
        RECT 115.970 111.305 116.140 111.845 ;
        RECT 111.280 110.920 112.880 111.090 ;
        RECT 114.310 110.920 115.910 111.090 ;
        RECT 78.560 110.680 80.160 110.850 ;
        RECT 81.590 110.680 83.190 110.850 ;
        RECT 97.230 110.720 98.830 110.890 ;
        RECT 100.260 110.720 101.860 110.890 ;
        RECT 64.510 110.480 66.110 110.650 ;
        RECT 67.540 110.480 69.140 110.650 ;
        RECT 103.790 107.170 105.390 107.340 ;
        RECT 106.820 107.170 108.420 107.340 ;
        RECT 71.070 106.930 72.670 107.100 ;
        RECT 74.100 106.930 75.700 107.100 ;
        RECT 70.840 106.075 71.010 106.715 ;
        RECT 72.730 106.075 72.900 106.715 ;
        RECT 73.870 106.075 74.040 106.715 ;
        RECT 75.760 106.075 75.930 106.715 ;
        RECT 103.560 106.315 103.730 106.955 ;
        RECT 105.450 106.315 105.620 106.955 ;
        RECT 106.590 106.315 106.760 106.955 ;
        RECT 108.480 106.315 108.650 106.955 ;
        RECT 103.790 105.930 105.390 106.100 ;
        RECT 106.820 105.930 108.420 106.100 ;
        RECT 71.070 105.690 72.670 105.860 ;
        RECT 74.100 105.690 75.700 105.860 ;
        RECT 103.190 102.860 104.790 103.030 ;
        RECT 106.220 102.860 107.820 103.030 ;
        RECT 70.470 102.620 72.070 102.790 ;
        RECT 70.240 101.210 70.410 102.450 ;
        RECT 72.130 101.210 72.300 102.450 ;
        RECT 73.270 101.210 73.440 102.450 ;
        RECT 75.160 101.210 75.330 102.450 ;
        RECT 102.960 101.450 103.130 102.690 ;
        RECT 104.850 101.450 105.020 102.690 ;
        RECT 105.990 101.450 106.160 102.690 ;
        RECT 107.880 101.450 108.050 102.690 ;
        RECT 103.190 101.110 104.790 101.280 ;
        RECT 106.220 101.110 107.820 101.280 ;
        RECT 70.470 100.870 72.070 101.040 ;
        RECT 98.040 97.330 99.640 97.500 ;
        RECT 101.070 97.330 102.670 97.500 ;
        RECT 65.320 97.090 66.920 97.260 ;
        RECT 68.350 97.090 69.950 97.260 ;
        RECT 65.090 96.460 65.260 96.920 ;
        RECT 70.010 96.460 70.180 96.920 ;
        RECT 97.810 96.700 97.980 97.160 ;
        RECT 102.730 96.700 102.900 97.160 ;
        RECT 98.040 96.360 99.640 96.530 ;
        RECT 101.070 96.360 102.670 96.530 ;
        RECT 65.320 96.120 66.920 96.290 ;
        RECT 68.350 96.120 69.950 96.290 ;
        RECT 109.930 85.960 111.530 86.130 ;
        RECT 112.960 85.960 114.560 86.130 ;
        RECT 95.880 85.760 97.480 85.930 ;
        RECT 98.910 85.760 100.510 85.930 ;
        RECT 95.650 85.005 95.820 85.545 ;
        RECT 100.570 85.005 100.740 85.545 ;
        RECT 109.700 85.205 109.870 85.745 ;
        RECT 114.620 85.205 114.790 85.745 ;
        RECT 109.930 84.820 111.530 84.990 ;
        RECT 112.960 84.820 114.560 84.990 ;
        RECT 95.880 84.620 97.480 84.790 ;
        RECT 98.910 84.620 100.510 84.790 ;
        RECT 78.280 83.440 79.880 83.610 ;
        RECT 81.310 83.440 82.910 83.610 ;
        RECT 64.230 83.240 65.830 83.410 ;
        RECT 67.260 83.240 68.860 83.410 ;
        RECT 64.000 82.485 64.170 83.025 ;
        RECT 68.920 82.485 69.090 83.025 ;
        RECT 78.050 82.685 78.220 83.225 ;
        RECT 82.970 82.685 83.140 83.225 ;
        RECT 78.280 82.300 79.880 82.470 ;
        RECT 81.310 82.300 82.910 82.470 ;
        RECT 64.230 82.100 65.830 82.270 ;
        RECT 67.260 82.100 68.860 82.270 ;
        RECT 102.440 81.070 104.040 81.240 ;
        RECT 105.470 81.070 107.070 81.240 ;
        RECT 102.210 80.215 102.380 80.855 ;
        RECT 104.100 80.215 104.270 80.855 ;
        RECT 105.240 80.215 105.410 80.855 ;
        RECT 107.130 80.215 107.300 80.855 ;
        RECT 102.440 79.830 104.040 80.000 ;
        RECT 105.470 79.830 107.070 80.000 ;
        RECT 70.790 78.550 72.390 78.720 ;
        RECT 73.820 78.550 75.420 78.720 ;
        RECT 70.560 77.695 70.730 78.335 ;
        RECT 72.450 77.695 72.620 78.335 ;
        RECT 73.590 77.695 73.760 78.335 ;
        RECT 75.480 77.695 75.650 78.335 ;
        RECT 70.790 77.310 72.390 77.480 ;
        RECT 73.820 77.310 75.420 77.480 ;
        RECT 101.840 76.760 103.440 76.930 ;
        RECT 104.870 76.760 106.470 76.930 ;
        RECT 101.610 75.350 101.780 76.590 ;
        RECT 103.500 75.350 103.670 76.590 ;
        RECT 104.640 75.350 104.810 76.590 ;
        RECT 106.530 75.350 106.700 76.590 ;
        RECT 101.840 75.010 103.440 75.180 ;
        RECT 104.870 75.010 106.470 75.180 ;
        RECT 70.190 74.240 71.790 74.410 ;
        RECT 69.960 72.830 70.130 74.070 ;
        RECT 71.850 72.830 72.020 74.070 ;
        RECT 72.990 72.830 73.160 74.070 ;
        RECT 74.880 72.830 75.050 74.070 ;
        RECT 70.190 72.490 71.790 72.660 ;
        RECT 96.690 71.230 98.290 71.400 ;
        RECT 99.720 71.230 101.320 71.400 ;
        RECT 96.460 70.600 96.630 71.060 ;
        RECT 101.380 70.600 101.550 71.060 ;
        RECT 96.690 70.260 98.290 70.430 ;
        RECT 99.720 70.260 101.320 70.430 ;
        RECT 65.040 68.710 66.640 68.880 ;
        RECT 68.070 68.710 69.670 68.880 ;
        RECT 64.810 68.080 64.980 68.540 ;
        RECT 69.730 68.080 69.900 68.540 ;
        RECT 65.040 67.740 66.640 67.910 ;
        RECT 68.070 67.740 69.670 67.910 ;
        RECT 72.570 58.970 74.170 59.140 ;
        RECT 75.600 58.970 77.200 59.140 ;
        RECT 72.340 58.260 72.510 58.800 ;
        RECT 74.230 58.260 74.400 58.800 ;
        RECT 75.370 58.260 75.540 58.800 ;
        RECT 77.260 58.260 77.430 58.800 ;
        RECT 72.570 57.920 74.170 58.090 ;
        RECT 75.600 57.920 77.200 58.090 ;
        RECT 86.980 57.810 88.580 57.980 ;
        RECT 90.010 57.810 91.610 57.980 ;
        RECT 86.750 57.100 86.920 57.640 ;
        RECT 88.640 57.100 88.810 57.640 ;
        RECT 89.780 57.100 89.950 57.640 ;
        RECT 91.670 57.100 91.840 57.640 ;
        RECT 72.570 56.900 74.170 57.070 ;
        RECT 75.600 56.900 77.200 57.070 ;
        RECT 86.980 56.760 88.580 56.930 ;
        RECT 90.010 56.760 91.610 56.930 ;
        RECT 72.340 56.190 72.510 56.730 ;
        RECT 77.260 56.190 77.430 56.730 ;
        RECT 72.570 55.850 74.170 56.020 ;
        RECT 75.600 55.850 77.200 56.020 ;
        RECT 86.980 55.740 88.580 55.910 ;
        RECT 90.010 55.740 91.610 55.910 ;
        RECT 86.750 55.030 86.920 55.570 ;
        RECT 91.670 55.030 91.840 55.570 ;
        RECT 86.980 54.690 88.580 54.860 ;
        RECT 90.010 54.690 91.610 54.860 ;
        RECT 80.750 43.170 82.350 43.340 ;
        RECT 83.780 43.170 85.380 43.340 ;
        RECT 80.520 42.415 80.690 42.955 ;
        RECT 85.440 42.415 85.610 42.955 ;
        RECT 80.750 42.030 82.350 42.200 ;
        RECT 83.780 42.030 85.380 42.200 ;
        RECT 80.750 41.010 82.350 41.180 ;
        RECT 83.780 41.010 85.380 41.180 ;
        RECT 80.520 40.255 80.690 40.795 ;
        RECT 85.440 40.255 85.610 40.795 ;
        RECT 80.750 39.870 82.350 40.040 ;
        RECT 83.780 39.870 85.380 40.040 ;
        RECT 77.980 34.380 89.280 34.550 ;
        RECT 77.980 19.120 78.150 34.380 ;
        RECT 89.110 19.120 89.280 34.380 ;
        RECT 77.980 18.950 89.280 19.120 ;
        RECT 89.750 34.450 101.050 34.620 ;
        RECT 89.750 19.190 89.920 34.450 ;
        RECT 100.880 19.190 101.050 34.450 ;
        RECT 89.750 19.020 101.050 19.190 ;
      LAYER met1 ;
        RECT 94.910 212.370 96.470 212.600 ;
        RECT 96.800 212.370 98.360 212.600 ;
        RECT 99.830 212.370 101.390 212.600 ;
        RECT 101.720 212.370 103.280 212.600 ;
        RECT 94.400 212.165 94.730 212.180 ;
        RECT 94.400 211.745 94.860 212.165 ;
        RECT 94.400 211.740 94.730 211.745 ;
        RECT 94.390 211.520 94.730 211.740 ;
        RECT 95.480 211.540 95.730 212.370 ;
        RECT 97.400 211.540 97.650 212.370 ;
        RECT 98.410 212.060 98.640 212.165 ;
        RECT 98.410 211.745 98.730 212.060 ;
        RECT 99.550 212.030 99.780 212.165 ;
        RECT 94.910 211.520 96.470 211.540 ;
        RECT 96.800 211.520 98.360 211.540 ;
        RECT 94.390 210.800 94.710 211.520 ;
        RECT 94.910 211.490 98.360 211.520 ;
        RECT 98.520 211.490 98.730 211.745 ;
        RECT 94.910 211.330 98.730 211.490 ;
        RECT 94.910 211.310 96.470 211.330 ;
        RECT 96.800 211.310 98.360 211.330 ;
        RECT 95.500 211.000 95.700 211.310 ;
        RECT 97.440 211.000 97.630 211.310 ;
        RECT 94.910 210.990 96.470 211.000 ;
        RECT 96.800 210.990 98.360 211.000 ;
        RECT 94.910 210.800 98.360 210.990 ;
        RECT 94.390 210.565 94.720 210.800 ;
        RECT 94.910 210.770 96.470 210.800 ;
        RECT 96.800 210.770 98.360 210.800 ;
        RECT 94.390 210.520 94.860 210.565 ;
        RECT 94.390 210.190 94.950 210.520 ;
        RECT 94.500 210.160 94.950 210.190 ;
        RECT 94.630 210.145 94.860 210.160 ;
        RECT 78.670 210.000 79.250 210.010 ;
        RECT 78.670 209.990 79.340 210.000 ;
        RECT 78.480 209.820 79.340 209.990 ;
        RECT 95.420 209.940 95.670 210.770 ;
        RECT 97.440 209.940 97.690 210.770 ;
        RECT 98.520 210.610 98.730 211.330 ;
        RECT 99.340 211.745 99.780 212.030 ;
        RECT 100.410 212.070 100.710 212.370 ;
        RECT 101.370 212.070 101.790 212.220 ;
        RECT 100.410 211.900 101.790 212.070 ;
        RECT 100.410 211.810 100.710 211.900 ;
        RECT 98.260 210.120 98.780 210.610 ;
        RECT 99.340 210.590 99.680 211.745 ;
        RECT 100.390 211.540 100.710 211.810 ;
        RECT 101.370 211.780 101.790 211.900 ;
        RECT 101.440 211.745 101.670 211.780 ;
        RECT 102.320 211.540 102.620 212.370 ;
        RECT 103.330 212.030 103.560 212.165 ;
        RECT 103.330 211.745 103.810 212.030 ;
        RECT 99.830 211.530 101.390 211.540 ;
        RECT 101.720 211.530 103.280 211.540 ;
        RECT 99.830 211.330 103.280 211.530 ;
        RECT 99.830 211.310 101.390 211.330 ;
        RECT 101.720 211.310 103.280 211.330 ;
        RECT 100.390 211.000 100.620 211.310 ;
        RECT 102.390 211.000 102.620 211.310 ;
        RECT 99.830 210.980 101.390 211.000 ;
        RECT 101.720 210.980 103.280 211.000 ;
        RECT 99.830 210.780 103.280 210.980 ;
        RECT 99.830 210.770 101.390 210.780 ;
        RECT 101.720 210.770 103.280 210.780 ;
        RECT 99.340 210.250 99.900 210.590 ;
        RECT 99.480 210.150 99.900 210.250 ;
        RECT 99.550 210.145 99.780 210.150 ;
        RECT 100.340 209.940 100.640 210.770 ;
        RECT 101.350 210.130 101.770 210.570 ;
        RECT 102.340 209.940 102.640 210.770 ;
        RECT 103.470 210.580 103.810 211.745 ;
        RECT 103.260 210.250 103.810 210.580 ;
        RECT 103.260 210.150 103.680 210.250 ;
        RECT 103.330 210.145 103.560 210.150 ;
        RECT 78.480 209.760 78.940 209.820 ;
        RECT 79.100 209.555 79.340 209.820 ;
        RECT 94.910 209.710 96.470 209.940 ;
        RECT 96.800 209.710 98.360 209.940 ;
        RECT 99.830 209.710 101.390 209.940 ;
        RECT 101.720 209.710 103.280 209.940 ;
        RECT 74.010 209.040 74.970 209.270 ;
        RECT 78.990 209.055 79.340 209.555 ;
        RECT 104.600 209.520 105.600 209.820 ;
        RECT 101.500 209.490 105.600 209.520 ;
        RECT 101.380 209.140 105.600 209.490 ;
        RECT 101.500 209.110 105.600 209.140 ;
        RECT 79.100 209.040 79.340 209.055 ;
        RECT 74.370 208.870 74.550 209.040 ;
        RECT 73.730 208.480 73.960 208.835 ;
        RECT 74.230 208.530 74.640 208.870 ;
        RECT 78.480 208.800 78.940 208.880 ;
        RECT 79.150 208.800 79.300 209.040 ;
        RECT 78.480 208.650 79.300 208.800 ;
        RECT 94.910 208.690 96.470 208.920 ;
        RECT 96.800 208.690 98.360 208.920 ;
        RECT 99.830 208.690 101.390 208.920 ;
        RECT 101.720 208.690 103.280 208.920 ;
        RECT 104.600 208.820 105.600 209.110 ;
        RECT 78.480 208.600 78.940 208.650 ;
        RECT 73.350 207.835 73.960 208.480 ;
        RECT 39.630 207.650 70.290 207.770 ;
        RECT 39.100 207.620 70.290 207.650 ;
        RECT 71.470 207.620 72.470 207.820 ;
        RECT 39.100 207.460 72.470 207.620 ;
        RECT 73.350 207.460 73.830 207.835 ;
        RECT 74.370 207.630 74.560 208.530 ;
        RECT 39.100 207.070 73.830 207.460 ;
        RECT 74.010 207.400 74.970 207.630 ;
        RECT 74.380 207.090 74.560 207.400 ;
        RECT 39.100 207.000 70.290 207.070 ;
        RECT 71.470 207.000 73.830 207.070 ;
        RECT 39.100 194.270 42.190 207.000 ;
        RECT 71.470 206.820 72.470 207.000 ;
        RECT 73.350 206.655 73.830 207.000 ;
        RECT 74.010 206.860 74.970 207.090 ;
        RECT 73.350 205.720 73.960 206.655 ;
        RECT 73.730 205.655 73.960 205.720 ;
        RECT 74.380 205.450 74.560 206.860 ;
        RECT 79.150 206.460 79.300 208.650 ;
        RECT 94.630 208.400 94.860 208.485 ;
        RECT 94.470 208.065 94.860 208.400 ;
        RECT 94.470 206.885 94.730 208.065 ;
        RECT 95.510 207.860 95.740 208.690 ;
        RECT 96.520 208.480 96.750 208.485 ;
        RECT 96.470 208.100 96.830 208.480 ;
        RECT 97.380 208.400 97.680 208.690 ;
        RECT 98.410 208.440 98.640 208.485 ;
        RECT 98.410 208.400 98.780 208.440 ;
        RECT 99.550 208.400 99.780 208.485 ;
        RECT 97.380 208.150 98.780 208.400 ;
        RECT 96.520 208.065 96.750 208.100 ;
        RECT 97.380 207.860 97.680 208.150 ;
        RECT 98.410 208.065 98.780 208.150 ;
        RECT 94.910 207.840 96.470 207.860 ;
        RECT 96.800 207.840 98.360 207.860 ;
        RECT 94.910 207.670 98.360 207.840 ;
        RECT 94.910 207.630 96.470 207.670 ;
        RECT 96.800 207.630 98.360 207.670 ;
        RECT 95.540 207.320 95.710 207.630 ;
        RECT 97.440 207.320 97.610 207.630 ;
        RECT 94.910 207.310 96.470 207.320 ;
        RECT 96.800 207.310 98.360 207.320 ;
        RECT 94.910 207.140 98.360 207.310 ;
        RECT 94.910 207.090 96.470 207.140 ;
        RECT 96.800 207.090 98.360 207.140 ;
        RECT 94.470 206.860 94.860 206.885 ;
        RECT 94.470 206.510 94.930 206.860 ;
        RECT 94.470 206.500 94.860 206.510 ;
        RECT 94.630 206.465 94.860 206.500 ;
        RECT 79.010 206.120 79.300 206.460 ;
        RECT 95.520 206.260 95.750 207.090 ;
        RECT 96.520 206.880 96.750 206.885 ;
        RECT 96.480 206.500 96.840 206.880 ;
        RECT 96.520 206.465 96.750 206.500 ;
        RECT 97.420 206.260 97.650 207.090 ;
        RECT 98.520 206.885 98.780 208.065 ;
        RECT 98.410 206.860 98.780 206.885 ;
        RECT 99.530 208.065 99.780 208.400 ;
        RECT 100.500 208.420 100.740 208.690 ;
        RECT 101.440 208.440 101.670 208.485 ;
        RECT 101.360 208.420 101.730 208.440 ;
        RECT 100.500 208.240 101.730 208.420 ;
        RECT 100.480 208.160 101.730 208.240 ;
        RECT 99.530 206.885 99.670 208.065 ;
        RECT 100.480 207.860 100.750 208.160 ;
        RECT 101.360 208.050 101.730 208.160 ;
        RECT 102.350 207.860 102.560 208.690 ;
        RECT 103.330 208.310 103.560 208.485 ;
        RECT 103.330 208.065 103.590 208.310 ;
        RECT 99.830 207.850 101.390 207.860 ;
        RECT 101.720 207.850 103.280 207.860 ;
        RECT 99.830 207.690 103.280 207.850 ;
        RECT 99.830 207.630 101.390 207.690 ;
        RECT 101.720 207.630 103.280 207.690 ;
        RECT 100.480 207.320 100.750 207.630 ;
        RECT 102.390 207.320 102.560 207.630 ;
        RECT 99.830 207.310 101.390 207.320 ;
        RECT 101.720 207.310 103.280 207.320 ;
        RECT 99.830 207.110 103.280 207.310 ;
        RECT 99.830 207.090 101.390 207.110 ;
        RECT 101.720 207.090 103.280 207.110 ;
        RECT 99.530 206.870 99.780 206.885 ;
        RECT 98.340 206.540 98.780 206.860 ;
        RECT 98.340 206.510 98.710 206.540 ;
        RECT 99.510 206.520 99.880 206.870 ;
        RECT 98.410 206.465 98.640 206.510 ;
        RECT 99.550 206.465 99.780 206.520 ;
        RECT 100.470 206.260 100.680 207.090 ;
        RECT 101.440 206.860 101.670 206.885 ;
        RECT 101.380 206.470 101.750 206.860 ;
        RECT 101.440 206.465 101.670 206.470 ;
        RECT 102.380 206.260 102.590 207.090 ;
        RECT 103.450 206.885 103.590 208.065 ;
        RECT 103.330 206.850 103.590 206.885 ;
        RECT 103.280 206.810 103.650 206.850 ;
        RECT 104.580 206.810 105.570 207.180 ;
        RECT 103.280 206.580 105.570 206.810 ;
        RECT 103.280 206.500 103.650 206.580 ;
        RECT 103.330 206.465 103.560 206.500 ;
        RECT 79.010 205.960 79.240 206.120 ;
        RECT 94.910 206.030 96.470 206.260 ;
        RECT 96.800 206.030 98.360 206.260 ;
        RECT 99.830 206.220 101.390 206.260 ;
        RECT 101.720 206.220 103.280 206.260 ;
        RECT 99.830 206.060 103.280 206.220 ;
        RECT 104.580 206.180 105.570 206.580 ;
        RECT 99.830 206.030 101.390 206.060 ;
        RECT 101.720 206.030 103.280 206.060 ;
        RECT 101.300 205.750 101.720 205.800 ;
        RECT 104.650 205.750 105.650 205.890 ;
        RECT 101.300 205.520 105.650 205.750 ;
        RECT 101.300 205.500 101.720 205.520 ;
        RECT 74.010 205.220 74.970 205.450 ;
        RECT 94.910 205.010 96.470 205.240 ;
        RECT 96.800 205.010 98.360 205.240 ;
        RECT 94.630 204.700 94.860 204.805 ;
        RECT 94.520 204.385 94.860 204.700 ;
        RECT 95.490 204.500 95.810 205.010 ;
        RECT 94.520 203.230 94.710 204.385 ;
        RECT 95.490 204.180 95.820 204.500 ;
        RECT 96.430 204.350 96.830 204.860 ;
        RECT 97.370 204.730 97.690 205.010 ;
        RECT 104.650 204.890 105.650 205.520 ;
        RECT 98.410 204.750 98.640 204.805 ;
        RECT 98.410 204.730 98.710 204.750 ;
        RECT 97.370 204.460 98.710 204.730 ;
        RECT 99.550 204.680 99.780 204.805 ;
        RECT 97.370 204.180 97.690 204.460 ;
        RECT 98.410 204.385 98.710 204.460 ;
        RECT 94.910 204.170 96.470 204.180 ;
        RECT 96.800 204.170 98.360 204.180 ;
        RECT 94.910 203.970 98.360 204.170 ;
        RECT 94.910 203.950 96.470 203.970 ;
        RECT 96.800 203.950 98.360 203.970 ;
        RECT 95.520 203.670 95.820 203.950 ;
        RECT 95.510 203.640 95.830 203.670 ;
        RECT 97.380 203.640 97.680 203.950 ;
        RECT 94.910 203.630 96.470 203.640 ;
        RECT 96.800 203.630 98.360 203.640 ;
        RECT 94.910 203.430 98.360 203.630 ;
        RECT 94.910 203.410 96.470 203.430 ;
        RECT 96.800 203.410 98.360 203.430 ;
        RECT 94.520 202.790 94.960 203.230 ;
        RECT 94.630 202.785 94.860 202.790 ;
        RECT 95.510 202.580 95.830 203.410 ;
        RECT 97.380 203.370 97.720 203.410 ;
        RECT 96.440 202.750 96.840 203.260 ;
        RECT 97.400 202.580 97.720 203.370 ;
        RECT 98.520 203.210 98.710 204.385 ;
        RECT 99.470 204.385 99.780 204.680 ;
        RECT 103.330 204.730 103.560 204.805 ;
        RECT 103.330 204.385 103.670 204.730 ;
        RECT 99.470 203.260 99.660 204.385 ;
        RECT 103.480 203.260 103.670 204.385 ;
        RECT 147.030 203.590 148.400 203.760 ;
        RECT 98.340 202.810 98.760 203.210 ;
        RECT 98.410 202.785 98.640 202.810 ;
        RECT 99.470 202.800 99.890 203.260 ;
        RECT 103.280 203.160 103.670 203.260 ;
        RECT 104.510 203.430 105.510 203.530 ;
        RECT 107.860 203.430 148.400 203.590 ;
        RECT 104.510 203.160 148.400 203.430 ;
        RECT 103.280 202.880 148.400 203.160 ;
        RECT 103.280 202.820 105.510 202.880 ;
        RECT 103.280 202.800 103.670 202.820 ;
        RECT 99.550 202.785 99.780 202.800 ;
        RECT 103.330 202.785 103.560 202.800 ;
        RECT 94.910 202.350 96.470 202.580 ;
        RECT 96.800 202.350 98.360 202.580 ;
        RECT 104.510 202.530 105.510 202.820 ;
        RECT 107.810 202.690 148.400 202.880 ;
        RECT 107.860 202.670 108.140 202.690 ;
        RECT 109.810 202.670 148.400 202.690 ;
        RECT 38.780 191.380 42.190 194.270 ;
        RECT 146.280 198.410 148.400 202.670 ;
        RECT 38.780 187.090 42.150 191.380 ;
        RECT 38.780 186.450 42.190 187.090 ;
        RECT 39.100 175.810 42.190 186.450 ;
        RECT 56.720 186.680 57.520 186.720 ;
        RECT 68.490 186.710 69.490 187.040 ;
        RECT 64.810 186.680 69.490 186.710 ;
        RECT 56.720 186.640 69.490 186.680 ;
        RECT 74.040 186.640 74.420 186.650 ;
        RECT 56.720 186.290 74.420 186.640 ;
        RECT 56.720 186.060 69.490 186.290 ;
        RECT 56.720 183.290 57.520 186.060 ;
        RECT 68.490 186.040 69.490 186.060 ;
        RECT 68.790 185.710 69.260 186.040 ;
        RECT 74.040 186.000 74.420 186.290 ;
        RECT 90.910 186.010 91.910 186.360 ;
        RECT 110.690 186.010 111.690 186.690 ;
        RECT 90.910 186.000 111.760 186.010 ;
        RECT 74.040 185.900 131.870 186.000 ;
        RECT 67.470 185.470 70.620 185.710 ;
        RECT 74.040 185.470 131.990 185.900 ;
        RECT 46.120 181.240 46.630 181.640 ;
        RECT 46.160 180.760 46.550 181.240 ;
        RECT 56.650 181.050 57.530 183.290 ;
        RECT 67.480 183.280 67.670 185.470 ;
        RECT 70.410 183.280 70.620 185.470 ;
        RECT 90.910 185.380 131.990 185.470 ;
        RECT 90.910 185.360 91.910 185.380 ;
        RECT 91.210 185.030 91.680 185.360 ;
        RECT 109.570 185.200 131.990 185.380 ;
        RECT 109.570 185.120 112.820 185.200 ;
        RECT 131.040 185.150 131.930 185.200 ;
        RECT 89.890 184.790 93.040 185.030 ;
        RECT 67.435 183.220 67.725 183.280 ;
        RECT 68.025 183.220 68.315 183.280 ;
        RECT 67.435 183.050 68.315 183.220 ;
        RECT 69.755 183.260 70.045 183.280 ;
        RECT 70.345 183.260 70.635 183.280 ;
        RECT 69.755 183.090 70.635 183.260 ;
        RECT 69.755 183.050 70.045 183.090 ;
        RECT 70.345 183.050 70.635 183.090 ;
        RECT 67.760 181.470 67.990 182.845 ;
        RECT 67.670 181.060 68.150 181.470 ;
        RECT 68.880 181.110 69.250 181.480 ;
        RECT 70.080 181.420 70.310 182.845 ;
        RECT 89.900 182.600 90.090 184.790 ;
        RECT 90.980 183.380 91.980 184.380 ;
        RECT 89.855 182.540 90.145 182.600 ;
        RECT 90.445 182.540 90.735 182.600 ;
        RECT 89.855 182.370 90.735 182.540 ;
        RECT 46.775 180.760 47.065 180.800 ;
        RECT 46.160 180.750 47.065 180.760 ;
        RECT 47.365 180.750 47.655 180.800 ;
        RECT 47.955 180.750 48.245 180.800 ;
        RECT 46.160 180.620 48.245 180.750 ;
        RECT 46.160 180.390 46.550 180.620 ;
        RECT 46.770 180.600 48.245 180.620 ;
        RECT 46.775 180.570 47.065 180.600 ;
        RECT 47.365 180.570 47.655 180.600 ;
        RECT 47.955 180.570 48.245 180.600 ;
        RECT 46.160 180.365 46.590 180.390 ;
        RECT 46.160 179.945 46.740 180.365 ;
        RECT 47.690 180.350 47.920 180.365 ;
        RECT 47.560 179.950 48.040 180.350 ;
        RECT 67.760 180.345 67.990 181.060 ;
        RECT 70.020 181.030 70.390 181.420 ;
        RECT 71.670 181.320 72.030 181.410 ;
        RECT 72.380 181.320 73.380 181.860 ;
        RECT 89.590 181.430 89.820 182.165 ;
        RECT 71.670 181.150 73.380 181.320 ;
        RECT 71.670 181.120 72.080 181.150 ;
        RECT 70.080 180.345 70.310 181.030 ;
        RECT 71.670 180.990 72.030 181.120 ;
        RECT 72.380 180.860 73.380 181.150 ;
        RECT 89.490 180.960 89.960 181.430 ;
        RECT 67.435 180.110 67.725 180.140 ;
        RECT 68.025 180.110 68.315 180.140 ;
        RECT 47.690 179.945 47.920 179.950 ;
        RECT 46.160 179.710 46.590 179.945 ;
        RECT 67.435 179.940 68.315 180.110 ;
        RECT 67.435 179.910 67.725 179.940 ;
        RECT 68.025 179.910 68.315 179.940 ;
        RECT 69.755 180.110 70.045 180.140 ;
        RECT 70.345 180.110 70.635 180.140 ;
        RECT 69.755 179.940 70.635 180.110 ;
        RECT 69.755 179.910 70.045 179.940 ;
        RECT 70.345 179.910 70.635 179.940 ;
        RECT 46.775 179.710 47.065 179.740 ;
        RECT 46.120 179.660 47.065 179.710 ;
        RECT 47.365 179.660 47.655 179.740 ;
        RECT 47.955 179.660 48.245 179.740 ;
        RECT 89.590 179.665 89.820 180.960 ;
        RECT 90.180 180.790 90.410 182.165 ;
        RECT 90.770 181.370 91.000 182.165 ;
        RECT 90.720 181.300 91.100 181.370 ;
        RECT 91.310 181.300 91.510 183.380 ;
        RECT 92.830 182.600 93.040 184.790 ;
        RECT 109.570 184.530 109.870 185.120 ;
        RECT 109.680 182.930 109.870 184.530 ;
        RECT 110.760 183.710 111.760 184.710 ;
        RECT 109.635 182.870 109.925 182.930 ;
        RECT 110.225 182.870 110.515 182.930 ;
        RECT 109.635 182.700 110.515 182.870 ;
        RECT 92.175 182.580 92.465 182.600 ;
        RECT 92.765 182.580 93.055 182.600 ;
        RECT 92.175 182.410 93.055 182.580 ;
        RECT 92.175 182.370 92.465 182.410 ;
        RECT 92.765 182.370 93.055 182.410 ;
        RECT 91.910 181.420 92.140 182.165 ;
        RECT 91.730 181.300 92.230 181.420 ;
        RECT 90.720 181.140 92.230 181.300 ;
        RECT 90.720 181.060 91.100 181.140 ;
        RECT 91.730 181.080 92.230 181.140 ;
        RECT 90.090 180.380 90.570 180.790 ;
        RECT 90.180 179.665 90.410 180.380 ;
        RECT 90.770 179.665 91.000 181.060 ;
        RECT 91.300 180.430 91.670 180.800 ;
        RECT 91.910 179.665 92.140 181.080 ;
        RECT 92.500 180.740 92.730 182.165 ;
        RECT 93.090 181.390 93.320 182.165 ;
        RECT 109.370 181.760 109.600 182.495 ;
        RECT 93.030 181.060 93.400 181.390 ;
        RECT 109.270 181.290 109.740 181.760 ;
        RECT 92.440 180.350 92.810 180.740 ;
        RECT 92.500 179.665 92.730 180.350 ;
        RECT 93.090 179.665 93.320 181.060 ;
        RECT 94.090 180.640 94.450 180.730 ;
        RECT 94.800 180.640 95.800 181.180 ;
        RECT 94.090 180.470 95.800 180.640 ;
        RECT 94.090 180.440 94.500 180.470 ;
        RECT 94.090 180.310 94.450 180.440 ;
        RECT 94.800 180.180 95.800 180.470 ;
        RECT 109.370 179.995 109.600 181.290 ;
        RECT 109.960 181.120 110.190 182.495 ;
        RECT 110.550 181.700 110.780 182.495 ;
        RECT 110.500 181.630 110.880 181.700 ;
        RECT 111.090 181.630 111.290 183.710 ;
        RECT 112.610 182.930 112.820 185.120 ;
        RECT 111.955 182.910 112.245 182.930 ;
        RECT 112.545 182.910 112.835 182.930 ;
        RECT 111.955 182.740 112.835 182.910 ;
        RECT 111.955 182.700 112.245 182.740 ;
        RECT 112.545 182.700 112.835 182.740 ;
        RECT 111.690 181.750 111.920 182.495 ;
        RECT 111.510 181.630 112.010 181.750 ;
        RECT 110.500 181.470 112.010 181.630 ;
        RECT 110.500 181.390 110.880 181.470 ;
        RECT 111.510 181.410 112.010 181.470 ;
        RECT 109.870 180.710 110.350 181.120 ;
        RECT 109.960 179.995 110.190 180.710 ;
        RECT 110.550 179.995 110.780 181.390 ;
        RECT 111.080 180.760 111.450 181.130 ;
        RECT 111.690 179.995 111.920 181.410 ;
        RECT 112.280 181.070 112.510 182.495 ;
        RECT 112.870 181.720 113.100 182.495 ;
        RECT 128.680 181.930 129.540 181.960 ;
        RECT 128.665 181.920 129.545 181.930 ;
        RECT 130.240 181.920 130.480 181.960 ;
        RECT 128.665 181.740 130.480 181.920 ;
        RECT 112.810 181.390 113.180 181.720 ;
        RECT 128.665 181.710 129.545 181.740 ;
        RECT 128.665 181.700 128.955 181.710 ;
        RECT 129.255 181.700 129.545 181.710 ;
        RECT 112.220 180.680 112.590 181.070 ;
        RECT 112.280 179.995 112.510 180.680 ;
        RECT 112.870 179.995 113.100 181.390 ;
        RECT 113.870 180.970 114.230 181.060 ;
        RECT 114.580 180.970 115.580 181.510 ;
        RECT 113.870 180.800 115.580 180.970 ;
        RECT 113.870 180.770 114.280 180.800 ;
        RECT 113.870 180.640 114.230 180.770 ;
        RECT 114.580 180.510 115.580 180.800 ;
        RECT 125.840 180.760 126.840 181.270 ;
        RECT 127.140 180.760 127.560 180.970 ;
        RECT 125.840 180.580 127.560 180.760 ;
        RECT 125.840 180.270 126.840 180.580 ;
        RECT 127.140 180.500 127.560 180.580 ;
        RECT 128.400 180.160 128.630 181.495 ;
        RECT 128.990 181.020 129.220 181.495 ;
        RECT 128.890 180.510 129.420 181.020 ;
        RECT 128.310 179.990 128.710 180.160 ;
        RECT 109.635 179.760 109.925 179.790 ;
        RECT 110.225 179.760 110.515 179.790 ;
        RECT 46.120 179.570 48.270 179.660 ;
        RECT 46.160 179.190 46.590 179.570 ;
        RECT 46.775 179.510 48.270 179.570 ;
        RECT 109.635 179.590 110.515 179.760 ;
        RECT 109.635 179.560 109.925 179.590 ;
        RECT 110.225 179.560 110.515 179.590 ;
        RECT 111.955 179.760 112.245 179.790 ;
        RECT 112.545 179.760 112.835 179.790 ;
        RECT 111.955 179.590 112.835 179.760 ;
        RECT 111.955 179.560 112.245 179.590 ;
        RECT 112.545 179.560 112.835 179.590 ;
        RECT 128.290 179.570 128.710 179.990 ;
        RECT 47.410 179.200 47.590 179.510 ;
        RECT 89.855 179.430 90.145 179.460 ;
        RECT 90.445 179.430 90.735 179.460 ;
        RECT 89.855 179.260 90.735 179.430 ;
        RECT 89.855 179.230 90.145 179.260 ;
        RECT 90.445 179.230 90.735 179.260 ;
        RECT 92.175 179.430 92.465 179.460 ;
        RECT 92.765 179.430 93.055 179.460 ;
        RECT 92.175 179.260 93.055 179.430 ;
        RECT 92.175 179.230 92.465 179.260 ;
        RECT 92.765 179.230 93.055 179.260 ;
        RECT 46.775 179.190 47.065 179.200 ;
        RECT 47.365 179.190 47.655 179.200 ;
        RECT 47.955 179.190 48.245 179.200 ;
        RECT 46.160 179.050 48.250 179.190 ;
        RECT 46.160 178.765 46.590 179.050 ;
        RECT 46.775 179.040 48.250 179.050 ;
        RECT 67.435 179.080 67.725 179.120 ;
        RECT 68.025 179.080 68.315 179.120 ;
        RECT 46.775 178.970 47.065 179.040 ;
        RECT 47.365 178.970 47.655 179.040 ;
        RECT 47.955 178.970 48.245 179.040 ;
        RECT 67.435 178.910 68.315 179.080 ;
        RECT 67.435 178.890 67.725 178.910 ;
        RECT 68.025 178.890 68.315 178.910 ;
        RECT 69.755 179.080 70.045 179.120 ;
        RECT 70.345 179.080 70.635 179.120 ;
        RECT 69.755 178.910 70.635 179.080 ;
        RECT 69.755 178.890 70.045 178.910 ;
        RECT 70.345 178.890 70.635 178.910 ;
        RECT 128.290 178.995 128.630 179.570 ;
        RECT 128.990 178.995 129.220 180.510 ;
        RECT 129.580 180.180 129.810 181.495 ;
        RECT 130.240 180.610 130.480 181.740 ;
        RECT 130.960 180.610 131.960 180.880 ;
        RECT 130.240 180.370 131.960 180.610 ;
        RECT 129.520 179.590 129.920 180.180 ;
        RECT 129.580 178.995 129.810 179.590 ;
        RECT 46.160 178.345 46.740 178.765 ;
        RECT 47.690 178.760 47.920 178.765 ;
        RECT 47.560 178.360 48.040 178.760 ;
        RECT 109.635 178.730 109.925 178.770 ;
        RECT 110.225 178.730 110.515 178.770 ;
        RECT 63.170 178.420 64.170 178.530 ;
        RECT 63.170 178.400 64.680 178.420 ;
        RECT 47.690 178.345 47.920 178.360 ;
        RECT 46.160 178.110 46.590 178.345 ;
        RECT 46.775 178.110 47.065 178.140 ;
        RECT 46.160 178.100 47.065 178.110 ;
        RECT 47.365 178.100 47.655 178.140 ;
        RECT 47.955 178.100 48.245 178.140 ;
        RECT 46.160 177.950 48.260 178.100 ;
        RECT 46.160 177.560 46.590 177.950 ;
        RECT 46.775 177.910 47.065 177.950 ;
        RECT 47.365 177.910 47.655 177.950 ;
        RECT 47.955 177.910 48.245 177.950 ;
        RECT 47.410 177.600 47.590 177.910 ;
        RECT 63.170 177.860 64.770 178.400 ;
        RECT 46.775 177.570 47.065 177.600 ;
        RECT 47.365 177.580 47.655 177.600 ;
        RECT 47.955 177.580 48.245 177.600 ;
        RECT 47.365 177.570 48.245 177.580 ;
        RECT 46.775 177.560 48.245 177.570 ;
        RECT 46.160 177.420 48.245 177.560 ;
        RECT 63.170 177.530 64.170 177.860 ;
        RECT 67.170 177.580 67.400 178.685 ;
        RECT 67.760 178.190 67.990 178.685 ;
        RECT 67.650 177.850 68.130 178.190 ;
        RECT 46.160 177.400 47.065 177.420 ;
        RECT 46.160 177.165 46.590 177.400 ;
        RECT 46.775 177.370 47.065 177.400 ;
        RECT 47.365 177.400 48.245 177.420 ;
        RECT 47.365 177.370 47.655 177.400 ;
        RECT 47.955 177.370 48.245 177.400 ;
        RECT 46.160 176.745 46.740 177.165 ;
        RECT 46.160 176.490 46.590 176.745 ;
        RECT 47.600 176.730 48.080 177.210 ;
        RECT 66.970 177.130 67.560 177.580 ;
        RECT 46.775 176.490 47.065 176.540 ;
        RECT 46.160 176.480 47.065 176.490 ;
        RECT 47.365 176.480 47.655 176.540 ;
        RECT 47.955 176.480 48.245 176.540 ;
        RECT 46.160 176.330 48.245 176.480 ;
        RECT 46.160 175.940 46.590 176.330 ;
        RECT 46.775 176.310 47.065 176.330 ;
        RECT 47.365 176.310 47.655 176.330 ;
        RECT 47.955 176.310 48.245 176.330 ;
        RECT 47.400 176.000 47.580 176.310 ;
        RECT 46.775 175.950 47.065 176.000 ;
        RECT 47.365 175.950 47.655 176.000 ;
        RECT 47.955 175.950 48.245 176.000 ;
        RECT 46.775 175.940 48.270 175.950 ;
        RECT 39.100 170.540 42.280 175.810 ;
        RECT 46.160 175.800 48.270 175.940 ;
        RECT 62.980 175.930 63.980 176.500 ;
        RECT 67.170 176.185 67.400 177.130 ;
        RECT 67.760 176.185 67.990 177.850 ;
        RECT 68.350 177.630 68.580 178.685 ;
        RECT 68.230 177.580 68.660 177.630 ;
        RECT 68.870 177.580 69.270 177.750 ;
        RECT 69.490 177.580 69.720 178.685 ;
        RECT 70.080 178.160 70.310 178.685 ;
        RECT 68.230 177.270 69.720 177.580 ;
        RECT 69.910 177.510 70.510 178.160 ;
        RECT 68.350 176.185 68.580 177.270 ;
        RECT 68.870 177.260 69.270 177.270 ;
        RECT 69.490 177.120 69.720 177.270 ;
        RECT 69.420 176.760 69.850 177.120 ;
        RECT 69.490 176.185 69.720 176.760 ;
        RECT 70.080 176.185 70.310 177.510 ;
        RECT 70.670 177.190 70.900 178.685 ;
        RECT 109.635 178.560 110.515 178.730 ;
        RECT 109.635 178.540 109.925 178.560 ;
        RECT 110.225 178.540 110.515 178.560 ;
        RECT 111.955 178.730 112.245 178.770 ;
        RECT 112.545 178.730 112.835 178.770 ;
        RECT 111.955 178.560 112.835 178.730 ;
        RECT 111.955 178.540 112.245 178.560 ;
        RECT 112.545 178.540 112.835 178.560 ;
        RECT 73.380 177.840 73.790 178.010 ;
        RECT 73.990 177.840 74.990 178.530 ;
        RECT 89.855 178.400 90.145 178.440 ;
        RECT 90.445 178.400 90.735 178.440 ;
        RECT 89.855 178.230 90.735 178.400 ;
        RECT 89.855 178.210 90.145 178.230 ;
        RECT 90.445 178.210 90.735 178.230 ;
        RECT 92.175 178.400 92.465 178.440 ;
        RECT 92.765 178.400 93.055 178.440 ;
        RECT 92.175 178.230 93.055 178.400 ;
        RECT 92.175 178.210 92.465 178.230 ;
        RECT 92.765 178.210 93.055 178.230 ;
        RECT 105.370 178.070 106.370 178.180 ;
        RECT 105.370 178.050 106.880 178.070 ;
        RECT 73.380 177.640 74.990 177.840 ;
        RECT 73.380 177.550 73.790 177.640 ;
        RECT 73.990 177.530 74.990 177.640 ;
        RECT 85.590 177.740 86.590 177.850 ;
        RECT 85.590 177.720 87.100 177.740 ;
        RECT 70.590 176.770 70.970 177.190 ;
        RECT 85.590 177.180 87.190 177.720 ;
        RECT 85.590 176.850 86.590 177.180 ;
        RECT 89.590 176.900 89.820 178.005 ;
        RECT 90.180 177.510 90.410 178.005 ;
        RECT 90.070 177.170 90.550 177.510 ;
        RECT 70.670 176.185 70.900 176.770 ;
        RECT 67.435 175.950 67.725 175.980 ;
        RECT 68.025 175.950 68.315 175.980 ;
        RECT 62.980 175.920 63.990 175.930 ;
        RECT 67.435 175.920 68.315 175.950 ;
        RECT 46.160 175.780 47.065 175.800 ;
        RECT 46.160 175.565 46.590 175.780 ;
        RECT 46.775 175.770 47.065 175.780 ;
        RECT 47.365 175.770 47.655 175.800 ;
        RECT 47.955 175.770 48.245 175.800 ;
        RECT 62.980 175.780 68.315 175.920 ;
        RECT 46.160 175.145 46.740 175.565 ;
        RECT 46.160 174.900 46.590 175.145 ;
        RECT 47.580 175.140 48.060 175.620 ;
        RECT 62.980 175.500 63.980 175.780 ;
        RECT 67.435 175.750 67.725 175.780 ;
        RECT 68.025 175.750 68.315 175.780 ;
        RECT 69.755 175.930 70.045 175.980 ;
        RECT 70.345 175.930 70.635 175.980 ;
        RECT 69.755 175.910 70.635 175.930 ;
        RECT 73.800 175.910 74.800 176.530 ;
        RECT 89.390 176.450 89.980 176.900 ;
        RECT 69.755 175.770 74.800 175.910 ;
        RECT 69.755 175.760 70.635 175.770 ;
        RECT 69.755 175.750 70.045 175.760 ;
        RECT 70.345 175.750 70.635 175.760 ;
        RECT 73.800 175.530 74.800 175.770 ;
        RECT 85.400 175.250 86.400 175.820 ;
        RECT 89.590 175.505 89.820 176.450 ;
        RECT 90.180 175.505 90.410 177.170 ;
        RECT 90.770 176.950 91.000 178.005 ;
        RECT 90.650 176.900 91.080 176.950 ;
        RECT 91.290 176.900 91.690 177.070 ;
        RECT 91.910 176.900 92.140 178.005 ;
        RECT 92.500 177.480 92.730 178.005 ;
        RECT 90.650 176.590 92.140 176.900 ;
        RECT 92.330 176.830 92.930 177.480 ;
        RECT 90.770 175.505 91.000 176.590 ;
        RECT 91.290 176.580 91.690 176.590 ;
        RECT 91.910 176.440 92.140 176.590 ;
        RECT 91.840 176.080 92.270 176.440 ;
        RECT 91.910 175.505 92.140 176.080 ;
        RECT 92.500 175.505 92.730 176.830 ;
        RECT 93.090 176.510 93.320 178.005 ;
        RECT 95.800 177.160 96.210 177.330 ;
        RECT 96.410 177.160 97.410 177.850 ;
        RECT 105.370 177.510 106.970 178.050 ;
        RECT 105.370 177.180 106.370 177.510 ;
        RECT 109.370 177.230 109.600 178.335 ;
        RECT 109.960 177.840 110.190 178.335 ;
        RECT 109.850 177.500 110.330 177.840 ;
        RECT 95.800 176.960 97.410 177.160 ;
        RECT 95.800 176.870 96.210 176.960 ;
        RECT 96.410 176.850 97.410 176.960 ;
        RECT 109.170 176.780 109.760 177.230 ;
        RECT 93.010 176.090 93.390 176.510 ;
        RECT 93.090 175.505 93.320 176.090 ;
        RECT 89.855 175.270 90.145 175.300 ;
        RECT 90.445 175.270 90.735 175.300 ;
        RECT 85.400 175.240 86.410 175.250 ;
        RECT 89.855 175.240 90.735 175.270 ;
        RECT 85.400 175.100 90.735 175.240 ;
        RECT 46.775 174.900 47.065 174.940 ;
        RECT 46.160 174.890 47.065 174.900 ;
        RECT 47.365 174.890 47.655 174.940 ;
        RECT 47.955 174.890 48.245 174.940 ;
        RECT 46.160 174.740 48.250 174.890 ;
        RECT 85.400 174.820 86.400 175.100 ;
        RECT 89.855 175.070 90.145 175.100 ;
        RECT 90.445 175.070 90.735 175.100 ;
        RECT 92.175 175.250 92.465 175.300 ;
        RECT 92.765 175.250 93.055 175.300 ;
        RECT 92.175 175.230 93.055 175.250 ;
        RECT 96.220 175.230 97.220 175.850 ;
        RECT 92.175 175.090 97.220 175.230 ;
        RECT 105.180 175.580 106.180 176.150 ;
        RECT 109.370 175.835 109.600 176.780 ;
        RECT 109.960 175.835 110.190 177.500 ;
        RECT 110.550 177.280 110.780 178.335 ;
        RECT 110.430 177.230 110.860 177.280 ;
        RECT 111.070 177.230 111.470 177.400 ;
        RECT 111.690 177.230 111.920 178.335 ;
        RECT 112.280 177.810 112.510 178.335 ;
        RECT 110.430 176.920 111.920 177.230 ;
        RECT 112.110 177.160 112.710 177.810 ;
        RECT 110.550 175.835 110.780 176.920 ;
        RECT 111.070 176.910 111.470 176.920 ;
        RECT 111.690 176.770 111.920 176.920 ;
        RECT 111.620 176.410 112.050 176.770 ;
        RECT 111.690 175.835 111.920 176.410 ;
        RECT 112.280 175.835 112.510 177.160 ;
        RECT 112.870 176.840 113.100 178.335 ;
        RECT 115.580 177.490 115.990 177.660 ;
        RECT 116.190 177.490 117.190 178.180 ;
        RECT 115.580 177.290 117.190 177.490 ;
        RECT 115.580 177.200 115.990 177.290 ;
        RECT 116.190 177.180 117.190 177.290 ;
        RECT 123.590 177.560 124.590 177.910 ;
        RECT 128.290 177.830 128.510 178.995 ;
        RECT 128.665 178.780 128.955 178.790 ;
        RECT 129.255 178.780 129.545 178.790 ;
        RECT 130.240 178.780 130.480 180.370 ;
        RECT 130.960 179.880 131.960 180.370 ;
        RECT 137.260 180.830 138.520 181.010 ;
        RECT 139.440 180.830 144.000 180.850 ;
        RECT 137.260 180.270 144.820 180.830 ;
        RECT 137.260 179.990 138.520 180.270 ;
        RECT 128.665 178.600 130.480 178.780 ;
        RECT 128.665 178.560 129.560 178.600 ;
        RECT 130.240 178.590 130.480 178.600 ;
        RECT 140.700 178.570 141.050 180.270 ;
        RECT 128.700 178.530 129.560 178.560 ;
        RECT 140.385 178.410 141.265 178.570 ;
        RECT 140.385 178.340 140.675 178.410 ;
        RECT 140.975 178.340 141.265 178.410 ;
        RECT 128.280 177.640 129.040 177.830 ;
        RECT 128.530 177.630 129.040 177.640 ;
        RECT 123.590 177.240 125.370 177.560 ;
        RECT 123.590 176.910 124.590 177.240 ;
        RECT 124.990 177.210 125.370 177.240 ;
        RECT 128.890 177.130 129.040 177.630 ;
        RECT 133.740 177.220 134.740 177.650 ;
        RECT 140.120 177.420 140.350 178.135 ;
        RECT 140.710 178.110 140.940 178.135 ;
        RECT 140.600 177.620 141.090 178.110 ;
        RECT 132.350 177.210 134.740 177.220 ;
        RECT 112.790 176.420 113.170 176.840 ;
        RECT 112.870 175.835 113.100 176.420 ;
        RECT 109.635 175.600 109.925 175.630 ;
        RECT 110.225 175.600 110.515 175.630 ;
        RECT 105.180 175.570 106.190 175.580 ;
        RECT 109.635 175.570 110.515 175.600 ;
        RECT 105.180 175.430 110.515 175.570 ;
        RECT 105.180 175.150 106.180 175.430 ;
        RECT 109.635 175.400 109.925 175.430 ;
        RECT 110.225 175.400 110.515 175.430 ;
        RECT 111.955 175.580 112.245 175.630 ;
        RECT 112.545 175.580 112.835 175.630 ;
        RECT 111.955 175.560 112.835 175.580 ;
        RECT 116.000 175.560 117.000 176.180 ;
        RECT 127.325 175.940 127.615 175.950 ;
        RECT 111.955 175.420 117.000 175.560 ;
        RECT 111.955 175.410 112.835 175.420 ;
        RECT 111.955 175.400 112.245 175.410 ;
        RECT 112.545 175.400 112.835 175.410 ;
        RECT 116.000 175.180 117.000 175.420 ;
        RECT 124.770 175.920 127.620 175.940 ;
        RECT 127.915 175.920 128.205 175.950 ;
        RECT 124.770 175.780 128.205 175.920 ;
        RECT 124.770 175.760 127.620 175.780 ;
        RECT 92.175 175.080 93.055 175.090 ;
        RECT 92.175 175.070 92.465 175.080 ;
        RECT 92.765 175.070 93.055 175.080 ;
        RECT 96.220 174.850 97.220 175.090 ;
        RECT 124.770 174.750 124.950 175.760 ;
        RECT 127.325 175.720 127.615 175.760 ;
        RECT 127.915 175.720 128.205 175.780 ;
        RECT 46.160 174.360 46.590 174.740 ;
        RECT 46.775 174.710 47.065 174.740 ;
        RECT 47.365 174.710 47.655 174.740 ;
        RECT 47.955 174.710 48.245 174.740 ;
        RECT 47.440 174.400 47.620 174.710 ;
        RECT 46.775 174.370 47.065 174.400 ;
        RECT 47.365 174.370 47.655 174.400 ;
        RECT 47.955 174.370 48.245 174.400 ;
        RECT 46.775 174.360 48.270 174.370 ;
        RECT 46.160 174.220 48.270 174.360 ;
        RECT 46.160 174.200 47.065 174.220 ;
        RECT 46.160 173.965 46.590 174.200 ;
        RECT 46.775 174.170 47.065 174.200 ;
        RECT 47.365 174.170 47.655 174.220 ;
        RECT 47.955 174.170 48.245 174.220 ;
        RECT 46.160 173.545 46.740 173.965 ;
        RECT 46.160 173.310 46.590 173.545 ;
        RECT 47.620 173.520 48.100 174.000 ;
        RECT 124.410 173.750 125.410 174.750 ;
        RECT 127.060 173.950 127.290 175.515 ;
        RECT 127.650 175.210 127.880 175.515 ;
        RECT 127.480 174.580 128.090 175.210 ;
        RECT 46.775 173.310 47.065 173.340 ;
        RECT 46.160 173.280 47.065 173.310 ;
        RECT 47.365 173.280 47.655 173.340 ;
        RECT 47.955 173.280 48.245 173.340 ;
        RECT 46.160 173.150 48.260 173.280 ;
        RECT 46.160 172.770 46.590 173.150 ;
        RECT 46.775 173.130 48.260 173.150 ;
        RECT 46.775 173.110 47.065 173.130 ;
        RECT 47.365 173.110 47.655 173.130 ;
        RECT 47.955 173.110 48.245 173.130 ;
        RECT 47.430 172.800 47.610 173.110 ;
        RECT 124.690 172.820 124.990 173.750 ;
        RECT 126.950 173.510 127.410 173.950 ;
        RECT 127.060 173.015 127.290 173.510 ;
        RECT 127.650 173.015 127.880 174.580 ;
        RECT 128.240 173.970 128.470 175.515 ;
        RECT 128.140 173.740 128.600 173.970 ;
        RECT 128.890 173.740 129.030 177.130 ;
        RECT 131.970 176.910 134.740 177.210 ;
        RECT 132.350 176.900 134.740 176.910 ;
        RECT 133.740 176.650 134.740 176.900 ;
        RECT 139.770 176.610 140.530 177.420 ;
        RECT 133.050 175.950 133.310 175.960 ;
        RECT 129.645 175.910 129.935 175.950 ;
        RECT 130.235 175.910 133.310 175.950 ;
        RECT 129.645 175.770 133.310 175.910 ;
        RECT 129.645 175.720 129.935 175.770 ;
        RECT 130.235 175.740 133.310 175.770 ;
        RECT 130.235 175.720 130.525 175.740 ;
        RECT 129.380 174.040 129.610 175.515 ;
        RECT 129.970 175.100 130.200 175.515 ;
        RECT 129.860 174.630 130.350 175.100 ;
        RECT 129.280 173.740 129.740 174.040 ;
        RECT 128.140 173.560 129.740 173.740 ;
        RECT 128.140 173.530 128.600 173.560 ;
        RECT 128.240 173.015 128.470 173.530 ;
        RECT 129.280 173.490 129.740 173.560 ;
        RECT 129.380 173.015 129.610 173.490 ;
        RECT 129.970 173.015 130.200 174.630 ;
        RECT 130.560 174.040 130.790 175.515 ;
        RECT 133.050 174.560 133.310 175.740 ;
        RECT 140.120 175.635 140.350 176.610 ;
        RECT 140.710 175.635 140.940 177.620 ;
        RECT 141.300 177.420 141.530 178.135 ;
        RECT 144.260 177.800 144.800 180.270 ;
        RECT 144.230 177.640 144.800 177.800 ;
        RECT 141.150 176.610 141.910 177.420 ;
        RECT 141.300 175.635 141.530 176.610 ;
        RECT 140.385 175.400 140.675 175.430 ;
        RECT 140.975 175.400 141.265 175.430 ;
        RECT 140.385 175.240 141.265 175.400 ;
        RECT 140.385 175.200 140.675 175.240 ;
        RECT 140.830 175.200 141.265 175.240 ;
        RECT 130.450 173.490 130.910 174.040 ;
        RECT 132.560 173.560 133.560 174.560 ;
        RECT 140.830 173.800 141.070 175.200 ;
        RECT 144.230 173.820 144.790 177.640 ;
        RECT 143.190 173.800 144.790 173.820 ;
        RECT 130.560 173.015 130.790 173.490 ;
        RECT 132.980 172.830 133.160 173.560 ;
        RECT 124.690 172.810 127.570 172.820 ;
        RECT 130.370 172.810 133.160 172.830 ;
        RECT 46.775 172.790 47.065 172.800 ;
        RECT 47.365 172.790 47.655 172.800 ;
        RECT 47.955 172.790 48.245 172.800 ;
        RECT 124.690 172.790 127.615 172.810 ;
        RECT 127.915 172.790 128.205 172.810 ;
        RECT 46.775 172.770 48.260 172.790 ;
        RECT 46.160 172.640 48.260 172.770 ;
        RECT 124.690 172.650 128.205 172.790 ;
        RECT 46.160 172.610 47.065 172.640 ;
        RECT 46.160 172.365 46.590 172.610 ;
        RECT 46.775 172.570 47.065 172.610 ;
        RECT 47.365 172.570 47.655 172.640 ;
        RECT 47.955 172.570 48.245 172.640 ;
        RECT 124.690 172.600 127.615 172.650 ;
        RECT 125.590 172.590 127.615 172.600 ;
        RECT 127.325 172.580 127.615 172.590 ;
        RECT 127.915 172.580 128.205 172.650 ;
        RECT 129.645 172.760 129.935 172.810 ;
        RECT 130.235 172.760 133.160 172.810 ;
        RECT 129.645 172.620 133.160 172.760 ;
        RECT 140.830 173.470 144.790 173.800 ;
        RECT 140.830 173.460 144.720 173.470 ;
        RECT 140.830 173.450 143.290 173.460 ;
        RECT 129.645 172.580 129.935 172.620 ;
        RECT 130.235 172.580 130.525 172.620 ;
        RECT 46.160 171.945 46.740 172.365 ;
        RECT 46.160 171.730 46.590 171.945 ;
        RECT 47.560 171.920 48.040 172.400 ;
        RECT 46.775 171.730 47.065 171.740 ;
        RECT 46.160 171.720 47.065 171.730 ;
        RECT 47.365 171.720 47.655 171.740 ;
        RECT 47.955 171.720 48.245 171.740 ;
        RECT 46.160 171.570 48.245 171.720 ;
        RECT 46.160 171.200 46.590 171.570 ;
        RECT 46.775 171.510 47.065 171.570 ;
        RECT 47.365 171.510 47.655 171.570 ;
        RECT 47.955 171.510 48.245 171.570 ;
        RECT 47.410 171.200 47.590 171.510 ;
        RECT 46.160 171.170 47.065 171.200 ;
        RECT 47.365 171.170 47.655 171.200 ;
        RECT 47.955 171.170 48.245 171.200 ;
        RECT 46.160 171.040 48.245 171.170 ;
        RECT 46.160 170.820 46.610 171.040 ;
        RECT 46.775 170.980 48.245 171.040 ;
        RECT 46.775 170.970 47.065 170.980 ;
        RECT 47.365 170.970 47.655 170.980 ;
        RECT 47.955 170.970 48.245 170.980 ;
        RECT 39.120 168.590 42.280 170.540 ;
        RECT 46.150 170.765 46.610 170.820 ;
        RECT 46.150 170.345 46.740 170.765 ;
        RECT 47.580 170.360 48.080 170.790 ;
        RECT 47.690 170.345 47.920 170.360 ;
        RECT 46.150 170.330 46.610 170.345 ;
        RECT 39.100 166.440 42.280 168.590 ;
        RECT 39.120 164.490 42.280 166.440 ;
        RECT 46.160 170.100 46.610 170.330 ;
        RECT 46.775 170.100 47.065 170.140 ;
        RECT 47.365 170.100 47.655 170.140 ;
        RECT 47.955 170.100 48.245 170.140 ;
        RECT 46.160 169.950 48.245 170.100 ;
        RECT 46.160 169.920 47.065 169.950 ;
        RECT 46.160 169.570 46.590 169.920 ;
        RECT 46.775 169.910 47.065 169.920 ;
        RECT 47.365 169.910 47.655 169.950 ;
        RECT 47.955 169.910 48.245 169.950 ;
        RECT 47.400 169.600 47.580 169.910 ;
        RECT 58.660 169.870 58.890 170.975 ;
        RECT 46.775 169.570 47.065 169.600 ;
        RECT 46.160 169.560 47.065 169.570 ;
        RECT 47.365 169.560 47.655 169.600 ;
        RECT 47.955 169.560 48.245 169.600 ;
        RECT 58.660 169.580 61.680 169.870 ;
        RECT 46.160 169.410 48.250 169.560 ;
        RECT 46.160 169.165 46.590 169.410 ;
        RECT 46.775 169.370 47.065 169.410 ;
        RECT 47.365 169.370 47.655 169.410 ;
        RECT 47.955 169.370 48.245 169.410 ;
        RECT 46.160 168.745 46.740 169.165 ;
        RECT 47.690 169.140 47.920 169.165 ;
        RECT 46.160 168.500 46.590 168.745 ;
        RECT 47.600 168.740 48.080 169.140 ;
        RECT 58.660 168.975 58.890 169.580 ;
        RECT 46.775 168.530 47.065 168.540 ;
        RECT 47.365 168.530 47.655 168.540 ;
        RECT 47.955 168.530 48.245 168.540 ;
        RECT 46.775 168.500 48.260 168.530 ;
        RECT 46.160 168.380 48.260 168.500 ;
        RECT 46.160 168.340 47.065 168.380 ;
        RECT 46.160 167.960 46.590 168.340 ;
        RECT 46.775 168.310 47.065 168.340 ;
        RECT 47.365 168.310 47.655 168.380 ;
        RECT 47.955 168.310 48.245 168.380 ;
        RECT 61.300 168.340 61.680 169.580 ;
        RECT 77.170 169.260 77.400 170.365 ;
        RECT 99.640 169.790 99.870 170.895 ;
        RECT 99.640 169.500 102.660 169.790 ;
        RECT 77.170 168.970 80.190 169.260 ;
        RECT 77.170 168.365 77.400 168.970 ;
        RECT 47.420 168.000 47.600 168.310 ;
        RECT 60.910 168.030 61.910 168.340 ;
        RECT 46.775 167.960 48.270 168.000 ;
        RECT 46.160 167.850 48.270 167.960 ;
        RECT 46.160 167.800 47.065 167.850 ;
        RECT 46.160 167.565 46.590 167.800 ;
        RECT 46.775 167.770 47.065 167.800 ;
        RECT 47.365 167.770 47.655 167.850 ;
        RECT 47.955 167.770 48.245 167.850 ;
        RECT 46.160 167.145 46.740 167.565 ;
        RECT 47.690 167.560 47.920 167.565 ;
        RECT 47.560 167.160 48.040 167.560 ;
        RECT 60.910 167.340 61.950 168.030 ;
        RECT 79.810 167.730 80.190 168.970 ;
        RECT 99.640 168.895 99.870 169.500 ;
        RECT 102.280 168.260 102.660 169.500 ;
        RECT 101.890 167.970 102.890 168.260 ;
        RECT 101.890 167.950 105.560 167.970 ;
        RECT 47.690 167.145 47.920 167.160 ;
        RECT 46.160 166.900 46.590 167.145 ;
        RECT 46.775 166.900 47.065 166.940 ;
        RECT 46.160 166.860 47.065 166.900 ;
        RECT 47.365 166.860 47.655 166.940 ;
        RECT 47.955 166.860 48.245 166.940 ;
        RECT 46.160 166.740 48.250 166.860 ;
        RECT 46.160 166.380 46.590 166.740 ;
        RECT 46.775 166.710 48.250 166.740 ;
        RECT 47.400 166.400 47.560 166.710 ;
        RECT 61.290 166.440 61.950 167.340 ;
        RECT 79.420 167.510 80.420 167.730 ;
        RECT 84.140 167.510 84.770 167.550 ;
        RECT 79.420 167.190 84.770 167.510 ;
        RECT 101.890 167.530 106.060 167.950 ;
        RECT 101.890 167.260 102.890 167.530 ;
        RECT 79.420 167.050 84.790 167.190 ;
        RECT 79.420 166.730 80.420 167.050 ;
        RECT 46.775 166.380 47.065 166.400 ;
        RECT 46.160 166.340 47.065 166.380 ;
        RECT 47.365 166.340 47.655 166.400 ;
        RECT 47.955 166.340 48.245 166.400 ;
        RECT 46.160 166.220 48.250 166.340 ;
        RECT 46.160 165.965 46.590 166.220 ;
        RECT 46.775 166.190 48.250 166.220 ;
        RECT 46.775 166.170 47.065 166.190 ;
        RECT 47.365 166.170 47.655 166.190 ;
        RECT 47.955 166.170 48.245 166.190 ;
        RECT 46.160 165.820 46.740 165.965 ;
        RECT 46.150 165.545 46.740 165.820 ;
        RECT 47.590 165.580 48.070 165.980 ;
        RECT 54.610 165.690 55.610 165.960 ;
        RECT 57.940 165.690 58.170 166.170 ;
        RECT 47.690 165.545 47.920 165.580 ;
        RECT 46.150 165.310 46.620 165.545 ;
        RECT 46.775 165.310 47.065 165.340 ;
        RECT 46.150 165.300 47.065 165.310 ;
        RECT 47.365 165.300 47.655 165.340 ;
        RECT 47.955 165.300 48.245 165.340 ;
        RECT 46.150 165.150 48.245 165.300 ;
        RECT 46.150 165.140 46.620 165.150 ;
        RECT 46.775 165.110 47.065 165.150 ;
        RECT 47.365 165.110 47.655 165.150 ;
        RECT 47.955 165.110 48.245 165.150 ;
        RECT 54.610 165.240 58.170 165.690 ;
        RECT 54.610 164.960 55.610 165.240 ;
        RECT 57.940 165.170 58.170 165.240 ;
        RECT 58.730 165.770 58.960 166.170 ;
        RECT 61.290 165.770 61.940 166.440 ;
        RECT 58.730 165.520 61.940 165.770 ;
        RECT 79.800 165.980 80.060 166.730 ;
        RECT 58.730 165.170 58.960 165.520 ;
        RECT 39.100 164.170 42.280 164.490 ;
        RECT 39.100 152.810 42.190 164.170 ;
        RECT 61.350 163.830 61.940 165.520 ;
        RECT 67.120 165.300 67.580 165.530 ;
        RECT 67.630 163.990 67.860 165.095 ;
        RECT 73.120 165.080 74.120 165.350 ;
        RECT 76.450 165.080 76.680 165.560 ;
        RECT 73.120 164.630 76.680 165.080 ;
        RECT 73.120 164.350 74.120 164.630 ;
        RECT 76.450 164.560 76.680 164.630 ;
        RECT 77.240 165.160 77.470 165.560 ;
        RECT 79.800 165.160 80.020 165.980 ;
        RECT 77.240 164.910 80.020 165.160 ;
        RECT 77.240 164.560 77.470 164.910 ;
        RECT 61.350 162.590 61.950 163.830 ;
        RECT 67.630 163.700 70.650 163.990 ;
        RECT 67.630 163.095 67.860 163.700 ;
        RECT 67.120 162.660 67.580 162.890 ;
        RECT 61.360 162.220 61.950 162.590 ;
        RECT 61.300 161.900 62.300 162.220 ;
        RECT 63.020 161.930 64.020 162.160 ;
        RECT 67.270 161.930 67.410 162.660 ;
        RECT 70.270 162.460 70.650 163.700 ;
        RECT 84.130 163.280 84.790 167.050 ;
        RECT 102.270 166.510 102.530 167.260 ;
        RECT 89.650 166.080 90.110 166.310 ;
        RECT 90.160 164.770 90.390 165.875 ;
        RECT 95.590 165.620 96.590 165.880 ;
        RECT 95.270 165.610 96.590 165.620 ;
        RECT 98.920 165.610 99.150 166.090 ;
        RECT 95.270 165.200 99.150 165.610 ;
        RECT 95.590 165.160 99.150 165.200 ;
        RECT 95.590 164.880 96.590 165.160 ;
        RECT 98.920 165.090 99.150 165.160 ;
        RECT 99.710 165.690 99.940 166.090 ;
        RECT 102.270 165.690 102.490 166.510 ;
        RECT 99.710 165.440 102.490 165.690 ;
        RECT 99.710 165.090 99.940 165.440 ;
        RECT 90.160 164.480 93.180 164.770 ;
        RECT 90.160 163.875 90.390 164.480 ;
        RECT 89.650 163.440 90.110 163.670 ;
        RECT 84.140 162.980 84.770 163.280 ;
        RECT 83.960 162.530 84.960 162.980 ;
        RECT 85.550 162.710 86.550 162.940 ;
        RECT 89.800 162.710 89.940 163.440 ;
        RECT 92.800 163.240 93.180 164.480 ;
        RECT 85.550 162.530 89.960 162.710 ;
        RECT 63.020 161.900 67.430 161.930 ;
        RECT 61.300 161.650 67.430 161.900 ;
        RECT 61.300 161.390 64.020 161.650 ;
        RECT 61.300 161.220 62.300 161.390 ;
        RECT 63.020 161.160 64.020 161.390 ;
        RECT 67.270 160.680 67.410 161.650 ;
        RECT 69.880 161.460 70.880 162.460 ;
        RECT 83.960 162.430 89.960 162.530 ;
        RECT 83.960 162.090 86.550 162.430 ;
        RECT 70.260 160.710 70.520 161.460 ;
        RECT 81.540 161.040 82.900 162.090 ;
        RECT 83.960 161.980 84.960 162.090 ;
        RECT 85.550 161.940 86.550 162.090 ;
        RECT 89.800 161.460 89.940 162.430 ;
        RECT 92.410 162.240 93.410 163.240 ;
        RECT 102.990 162.270 104.120 163.490 ;
        RECT 105.440 163.080 106.060 167.530 ;
        RECT 140.830 167.510 141.070 173.450 ;
        RECT 140.810 167.280 143.980 167.510 ;
        RECT 110.590 166.570 111.050 166.800 ;
        RECT 111.100 165.260 111.330 166.365 ;
        RECT 128.020 166.240 128.480 166.470 ;
        RECT 111.100 164.970 114.120 165.260 ;
        RECT 111.100 164.365 111.330 164.970 ;
        RECT 110.590 163.930 111.050 164.160 ;
        RECT 106.490 163.380 107.490 163.430 ;
        RECT 106.480 163.200 107.490 163.380 ;
        RECT 110.740 163.200 110.880 163.930 ;
        RECT 113.740 163.730 114.120 164.970 ;
        RECT 128.530 164.930 128.760 166.035 ;
        RECT 140.830 165.830 141.070 167.280 ;
        RECT 140.830 165.790 141.125 165.830 ;
        RECT 141.425 165.790 141.715 165.830 ;
        RECT 140.830 165.740 141.715 165.790 ;
        RECT 140.835 165.630 141.715 165.740 ;
        RECT 140.835 165.600 141.125 165.630 ;
        RECT 141.425 165.600 141.715 165.630 ;
        RECT 140.570 165.200 140.800 165.395 ;
        RECT 128.530 164.640 131.550 164.930 ;
        RECT 128.530 164.035 128.760 164.640 ;
        RECT 106.480 163.080 110.900 163.200 ;
        RECT 105.390 162.920 110.900 163.080 ;
        RECT 105.390 162.630 107.490 162.920 ;
        RECT 92.790 161.490 93.050 162.240 ;
        RECT 89.720 161.230 90.180 161.460 ;
        RECT 67.190 160.450 67.650 160.680 ;
        RECT 46.570 159.940 46.800 160.130 ;
        RECT 46.410 159.870 46.940 159.940 ;
        RECT 46.100 159.460 46.940 159.870 ;
        RECT 46.100 158.460 46.800 159.460 ;
        RECT 47.160 159.140 47.390 160.130 ;
        RECT 47.750 159.980 47.980 160.130 ;
        RECT 47.580 159.500 48.110 159.980 ;
        RECT 46.990 158.660 47.520 159.140 ;
        RECT 47.160 158.460 47.390 158.660 ;
        RECT 47.750 158.460 47.980 159.500 ;
        RECT 48.340 159.140 48.570 160.130 ;
        RECT 63.580 159.810 64.580 160.080 ;
        RECT 66.910 159.810 67.140 160.290 ;
        RECT 63.580 159.360 67.140 159.810 ;
        RECT 48.180 158.660 48.710 159.140 ;
        RECT 63.580 159.080 64.580 159.360 ;
        RECT 66.910 159.290 67.140 159.360 ;
        RECT 67.700 159.890 67.930 160.290 ;
        RECT 70.260 159.890 70.480 160.710 ;
        RECT 67.700 159.640 70.480 159.890 ;
        RECT 67.700 159.290 67.930 159.640 ;
        RECT 81.540 159.560 82.950 161.040 ;
        RECT 86.110 160.590 87.110 160.860 ;
        RECT 89.440 160.590 89.670 161.070 ;
        RECT 86.110 160.140 89.670 160.590 ;
        RECT 86.110 159.860 87.110 160.140 ;
        RECT 48.340 158.460 48.570 158.660 ;
        RECT 46.100 158.250 46.600 158.460 ;
        RECT 46.020 157.770 46.600 158.250 ;
        RECT 46.100 157.370 46.600 157.770 ;
        RECT 46.100 157.190 46.800 157.370 ;
        RECT 46.100 156.790 46.940 157.190 ;
        RECT 46.100 156.740 46.800 156.790 ;
        RECT 46.570 155.700 46.800 156.740 ;
        RECT 47.160 156.380 47.390 157.370 ;
        RECT 47.750 157.250 47.980 157.370 ;
        RECT 47.650 156.850 48.160 157.250 ;
        RECT 47.060 155.980 47.570 156.380 ;
        RECT 47.160 155.700 47.390 155.980 ;
        RECT 47.750 155.700 47.980 156.850 ;
        RECT 48.340 156.380 48.570 157.370 ;
        RECT 48.340 156.330 48.860 156.380 ;
        RECT 48.240 155.930 48.860 156.330 ;
        RECT 48.340 155.700 48.860 155.930 ;
        RECT 48.500 153.870 48.860 155.700 ;
        RECT 63.630 155.390 64.400 159.080 ;
        RECT 67.190 158.900 67.650 159.130 ;
        RECT 48.350 153.660 49.350 153.870 ;
        RECT 63.550 153.660 64.410 155.390 ;
        RECT 48.350 153.050 64.410 153.660 ;
        RECT 81.540 153.080 82.900 159.560 ;
        RECT 87.840 156.450 88.380 160.140 ;
        RECT 89.440 160.070 89.670 160.140 ;
        RECT 90.230 160.670 90.460 161.070 ;
        RECT 92.790 160.670 93.010 161.490 ;
        RECT 90.230 160.420 93.010 160.670 ;
        RECT 90.230 160.070 90.460 160.420 ;
        RECT 89.720 159.680 90.180 159.910 ;
        RECT 103.290 158.900 103.920 162.270 ;
        RECT 105.460 160.960 105.920 162.630 ;
        RECT 106.490 162.430 107.490 162.630 ;
        RECT 110.740 161.950 110.880 162.920 ;
        RECT 113.350 162.730 114.350 163.730 ;
        RECT 128.020 163.600 128.480 163.830 ;
        RECT 123.920 162.900 124.920 163.100 ;
        RECT 123.210 162.870 124.920 162.900 ;
        RECT 128.170 162.870 128.310 163.600 ;
        RECT 131.170 163.400 131.550 164.640 ;
        RECT 140.300 164.550 140.950 165.200 ;
        RECT 123.210 162.840 128.330 162.870 ;
        RECT 113.730 161.980 113.990 162.730 ;
        RECT 123.030 162.590 128.330 162.840 ;
        RECT 123.030 162.490 124.920 162.590 ;
        RECT 110.660 161.720 111.120 161.950 ;
        RECT 107.050 161.080 108.050 161.350 ;
        RECT 110.380 161.080 110.610 161.560 ;
        RECT 105.240 159.960 106.240 160.960 ;
        RECT 107.050 160.630 110.610 161.080 ;
        RECT 107.050 160.350 108.050 160.630 ;
        RECT 110.380 160.560 110.610 160.630 ;
        RECT 111.170 161.160 111.400 161.560 ;
        RECT 113.730 161.160 113.950 161.980 ;
        RECT 111.170 160.910 113.950 161.160 ;
        RECT 123.030 161.100 123.370 162.490 ;
        RECT 123.920 162.100 124.920 162.490 ;
        RECT 128.170 161.620 128.310 162.590 ;
        RECT 130.780 162.400 131.780 163.400 ;
        RECT 140.570 162.895 140.800 164.550 ;
        RECT 141.160 163.750 141.390 165.395 ;
        RECT 141.750 165.320 141.980 165.395 ;
        RECT 141.610 164.670 142.260 165.320 ;
        RECT 141.060 163.320 141.450 163.750 ;
        RECT 141.160 162.895 141.390 163.320 ;
        RECT 141.750 162.895 141.980 164.670 ;
        RECT 143.520 163.440 143.960 167.280 ;
        RECT 140.835 162.650 141.125 162.690 ;
        RECT 141.425 162.660 141.715 162.690 ;
        RECT 143.520 162.660 143.920 163.440 ;
        RECT 141.425 162.650 143.920 162.660 ;
        RECT 140.835 162.490 143.920 162.650 ;
        RECT 140.835 162.460 141.125 162.490 ;
        RECT 141.425 162.460 143.920 162.490 ;
        RECT 141.460 162.430 143.920 162.460 ;
        RECT 131.160 161.650 131.420 162.400 ;
        RECT 128.090 161.390 128.550 161.620 ;
        RECT 111.170 160.560 111.400 160.910 ;
        RECT 122.750 160.870 123.750 161.100 ;
        RECT 119.990 160.660 123.750 160.870 ;
        RECT 97.700 158.740 103.920 158.900 ;
        RECT 97.650 158.350 103.920 158.740 ;
        RECT 97.650 158.100 103.890 158.350 ;
        RECT 87.840 155.780 88.510 156.450 ;
        RECT 48.350 152.870 49.350 153.050 ;
        RECT 39.100 151.780 42.150 152.810 ;
        RECT 38.990 143.210 42.150 151.780 ;
        RECT 63.550 148.590 64.410 153.050 ;
        RECT 81.430 152.090 82.900 153.080 ;
        RECT 81.430 151.600 82.760 152.090 ;
        RECT 87.880 148.910 88.510 155.780 ;
        RECT 97.650 153.580 98.290 158.100 ;
        RECT 107.070 154.800 107.930 160.350 ;
        RECT 110.660 160.170 111.120 160.400 ;
        RECT 119.970 160.390 123.750 160.660 ;
        RECT 119.970 158.060 120.370 160.390 ;
        RECT 122.750 160.100 123.750 160.390 ;
        RECT 124.480 160.750 125.480 161.020 ;
        RECT 127.810 160.750 128.040 161.230 ;
        RECT 124.480 160.300 128.040 160.750 ;
        RECT 124.480 160.020 125.480 160.300 ;
        RECT 127.810 160.230 128.040 160.300 ;
        RECT 128.600 160.830 128.830 161.230 ;
        RECT 131.160 160.830 131.380 161.650 ;
        RECT 128.600 160.580 131.380 160.830 ;
        RECT 128.600 160.230 128.830 160.580 ;
        RECT 115.220 156.810 115.450 157.915 ;
        RECT 119.940 157.750 120.370 158.060 ;
        RECT 115.220 156.520 118.240 156.810 ;
        RECT 115.220 155.915 115.450 156.520 ;
        RECT 117.860 155.280 118.240 156.520 ;
        RECT 107.040 153.810 107.930 154.800 ;
        RECT 117.470 154.940 118.470 155.280 ;
        RECT 119.940 154.940 120.310 157.750 ;
        RECT 121.120 155.860 122.360 157.390 ;
        RECT 117.470 154.500 120.310 154.940 ;
        RECT 117.470 154.440 119.710 154.500 ;
        RECT 117.470 154.280 118.470 154.440 ;
        RECT 97.610 153.350 98.510 153.580 ;
        RECT 93.110 152.850 94.110 153.180 ;
        RECT 97.370 152.850 98.610 153.350 ;
        RECT 101.700 153.340 102.600 153.460 ;
        RECT 93.110 152.630 98.610 152.850 ;
        RECT 93.110 152.180 94.110 152.630 ;
        RECT 97.370 151.690 98.610 152.630 ;
        RECT 101.500 152.820 102.740 153.340 ;
        RECT 104.280 152.820 105.280 153.060 ;
        RECT 101.500 152.170 105.280 152.820 ;
        RECT 107.040 152.700 107.920 153.810 ;
        RECT 117.850 153.530 118.110 154.280 ;
        RECT 107.040 152.330 107.930 152.700 ;
        RECT 97.610 151.475 98.510 151.690 ;
        RECT 101.500 151.680 102.740 152.170 ;
        RECT 104.280 152.060 105.280 152.170 ;
        RECT 101.700 151.355 102.600 151.680 ;
        RECT 97.610 148.910 98.510 149.775 ;
        RECT 101.700 148.910 102.600 149.655 ;
        RECT 81.310 148.890 103.300 148.910 ;
        RECT 107.070 148.890 107.930 152.330 ;
        RECT 111.170 152.630 112.170 152.900 ;
        RECT 114.500 152.630 114.730 153.110 ;
        RECT 111.170 152.180 114.730 152.630 ;
        RECT 111.170 151.900 112.170 152.180 ;
        RECT 114.500 152.110 114.730 152.180 ;
        RECT 115.290 152.710 115.520 153.110 ;
        RECT 117.850 152.710 118.070 153.530 ;
        RECT 115.290 152.460 118.070 152.710 ;
        RECT 115.290 152.110 115.520 152.460 ;
        RECT 111.320 148.890 112.100 151.900 ;
        RECT 121.520 150.930 122.010 155.860 ;
        RECT 121.270 149.940 122.610 150.930 ;
        RECT 124.570 149.390 125.430 160.020 ;
        RECT 128.090 159.840 128.550 160.070 ;
        RECT 130.350 150.960 131.750 153.050 ;
        RECT 124.570 149.060 125.390 149.390 ;
        RECT 124.190 148.950 125.390 149.060 ;
        RECT 123.740 148.890 125.390 148.950 ;
        RECT 81.310 148.590 125.390 148.890 ;
        RECT 63.550 147.450 125.390 148.590 ;
        RECT 63.550 147.360 103.300 147.450 ;
        RECT 123.740 147.420 125.390 147.450 ;
        RECT 63.550 147.330 85.690 147.360 ;
        RECT 124.190 147.350 125.390 147.420 ;
        RECT 63.550 147.300 64.410 147.330 ;
        RECT 39.100 138.040 42.150 143.210 ;
        RECT 60.350 142.470 71.400 142.540 ;
        RECT 60.190 142.390 71.400 142.470 ;
        RECT 93.140 142.390 95.030 142.550 ;
        RECT 60.190 140.430 95.030 142.390 ;
        RECT 130.400 141.440 131.520 150.960 ;
        RECT 146.280 142.510 148.210 198.410 ;
        RECT 146.280 141.780 148.190 142.510 ;
        RECT 130.120 141.080 132.010 141.440 ;
        RECT 60.190 140.110 71.400 140.430 ;
        RECT 39.100 100.100 42.190 138.040 ;
        RECT 56.630 102.830 58.800 104.900 ;
        RECT 60.190 102.830 62.550 140.110 ;
        RECT 93.140 139.950 95.030 140.430 ;
        RECT 130.050 140.270 132.010 141.080 ;
        RECT 130.120 139.530 132.010 140.270 ;
        RECT 130.330 137.430 131.810 139.530 ;
        RECT 136.430 137.860 148.270 141.780 ;
        RECT 95.450 136.210 131.810 137.430 ;
        RECT 95.510 125.770 96.200 136.210 ;
        RECT 130.330 136.040 131.810 136.210 ;
        RECT 95.540 122.550 96.170 125.770 ;
        RECT 95.540 121.940 96.190 122.550 ;
        RECT 71.850 113.150 75.710 113.190 ;
        RECT 71.850 112.910 79.530 113.150 ;
        RECT 68.040 112.610 68.640 112.910 ;
        RECT 68.190 111.820 68.430 112.610 ;
        RECT 64.530 111.590 66.090 111.820 ;
        RECT 67.560 111.590 69.120 111.820 ;
        RECT 64.250 111.380 64.480 111.385 ;
        RECT 64.030 110.885 64.480 111.380 ;
        RECT 64.030 109.790 64.350 110.885 ;
        RECT 65.190 110.830 65.390 111.590 ;
        RECT 68.190 111.500 68.430 111.590 ;
        RECT 65.190 110.680 65.400 110.830 ;
        RECT 68.210 110.750 68.410 111.500 ;
        RECT 69.170 111.380 69.400 111.385 ;
        RECT 69.170 110.885 69.520 111.380 ;
        RECT 68.180 110.680 68.410 110.750 ;
        RECT 64.530 110.450 66.090 110.680 ;
        RECT 67.560 110.450 69.120 110.680 ;
        RECT 65.200 109.790 65.400 110.450 ;
        RECT 64.030 109.750 65.400 109.790 ;
        RECT 68.180 109.750 68.380 110.450 ;
        RECT 64.030 109.520 68.380 109.750 ;
        RECT 64.030 109.500 68.360 109.520 ;
        RECT 64.030 108.300 64.350 109.500 ;
        RECT 65.200 109.490 68.360 109.500 ;
        RECT 69.290 109.370 69.520 110.885 ;
        RECT 69.270 109.150 70.980 109.370 ;
        RECT 70.700 108.870 70.980 109.150 ;
        RECT 64.020 104.560 64.360 108.300 ;
        RECT 70.720 106.910 70.950 108.870 ;
        RECT 71.850 107.740 72.130 112.910 ;
        RECT 75.630 112.890 79.530 112.910 ;
        RECT 79.270 112.020 79.490 112.890 ;
        RECT 74.630 111.470 75.340 112.000 ;
        RECT 78.580 111.790 80.140 112.020 ;
        RECT 81.610 111.790 83.170 112.020 ;
        RECT 79.270 111.640 79.490 111.790 ;
        RECT 78.130 111.585 78.420 111.630 ;
        RECT 71.860 107.330 72.100 107.740 ;
        RECT 71.850 107.130 72.110 107.330 ;
        RECT 74.780 107.130 75.060 111.470 ;
        RECT 78.130 111.085 78.530 111.585 ;
        RECT 78.130 109.900 78.420 111.085 ;
        RECT 79.280 110.920 79.480 111.640 ;
        RECT 79.260 110.880 79.520 110.920 ;
        RECT 82.280 110.880 82.480 111.790 ;
        RECT 83.220 111.510 83.450 111.585 ;
        RECT 83.220 111.085 83.620 111.510 ;
        RECT 78.580 110.650 80.140 110.880 ;
        RECT 81.610 110.650 83.170 110.880 ;
        RECT 79.260 110.290 79.520 110.650 ;
        RECT 82.320 110.290 82.460 110.650 ;
        RECT 79.260 110.230 82.480 110.290 ;
        RECT 83.350 110.230 83.620 111.085 ;
        RECT 79.260 110.000 83.620 110.230 ;
        RECT 82.470 109.940 83.620 110.000 ;
        RECT 78.130 109.730 78.400 109.900 ;
        RECT 75.860 109.450 78.400 109.730 ;
        RECT 75.860 107.580 76.180 109.450 ;
        RECT 83.350 108.950 83.620 109.940 ;
        RECT 83.350 108.430 83.640 108.950 ;
        RECT 70.730 106.695 70.940 106.910 ;
        RECT 71.090 106.900 72.650 107.130 ;
        RECT 74.120 106.900 75.680 107.130 ;
        RECT 70.730 106.240 71.040 106.695 ;
        RECT 70.810 106.095 71.040 106.240 ;
        RECT 71.850 105.890 72.110 106.900 ;
        RECT 72.700 106.510 72.930 106.695 ;
        RECT 73.840 106.510 74.070 106.695 ;
        RECT 72.700 106.330 74.070 106.510 ;
        RECT 72.700 106.095 72.930 106.330 ;
        RECT 71.090 105.660 72.650 105.890 ;
        RECT 73.220 104.900 73.490 106.330 ;
        RECT 73.840 106.095 74.070 106.330 ;
        RECT 74.770 105.890 75.090 106.900 ;
        RECT 75.870 106.695 76.180 107.580 ;
        RECT 75.730 106.180 76.180 106.695 ;
        RECT 75.730 106.095 75.960 106.180 ;
        RECT 83.370 106.020 83.640 108.430 ;
        RECT 95.630 107.170 96.190 121.940 ;
        RECT 104.570 113.390 108.430 113.430 ;
        RECT 104.570 113.150 112.250 113.390 ;
        RECT 100.760 112.850 101.360 113.150 ;
        RECT 100.910 112.060 101.150 112.850 ;
        RECT 97.250 111.830 98.810 112.060 ;
        RECT 100.280 111.830 101.840 112.060 ;
        RECT 96.970 111.620 97.200 111.625 ;
        RECT 96.750 111.125 97.200 111.620 ;
        RECT 96.750 110.030 97.070 111.125 ;
        RECT 97.910 111.070 98.110 111.830 ;
        RECT 100.910 111.740 101.150 111.830 ;
        RECT 97.910 110.920 98.120 111.070 ;
        RECT 100.930 110.990 101.130 111.740 ;
        RECT 101.890 111.620 102.120 111.625 ;
        RECT 101.890 111.125 102.240 111.620 ;
        RECT 100.900 110.920 101.130 110.990 ;
        RECT 97.250 110.690 98.810 110.920 ;
        RECT 100.280 110.690 101.840 110.920 ;
        RECT 97.920 110.030 98.120 110.690 ;
        RECT 96.750 109.990 98.120 110.030 ;
        RECT 100.900 109.990 101.100 110.690 ;
        RECT 96.750 109.760 101.100 109.990 ;
        RECT 96.750 109.740 101.080 109.760 ;
        RECT 96.750 108.540 97.070 109.740 ;
        RECT 97.920 109.730 101.080 109.740 ;
        RECT 102.010 109.610 102.240 111.125 ;
        RECT 101.990 109.390 103.700 109.610 ;
        RECT 103.420 109.110 103.700 109.390 ;
        RECT 88.780 106.460 96.200 107.170 ;
        RECT 74.120 105.660 75.680 105.890 ;
        RECT 64.040 104.220 64.360 104.560 ;
        RECT 64.040 104.080 70.300 104.220 ;
        RECT 64.040 104.010 70.310 104.080 ;
        RECT 64.040 104.000 64.360 104.010 ;
        RECT 56.630 102.810 64.490 102.830 ;
        RECT 67.890 102.810 68.890 102.910 ;
        RECT 56.630 102.230 68.890 102.810 ;
        RECT 56.630 102.000 58.800 102.230 ;
        RECT 60.190 102.160 68.890 102.230 ;
        RECT 67.890 101.910 68.890 102.160 ;
        RECT 70.130 102.430 70.310 104.010 ;
        RECT 72.920 103.900 73.920 104.900 ;
        RECT 83.370 103.740 83.650 106.020 ;
        RECT 75.250 103.590 83.650 103.740 ;
        RECT 75.240 103.460 83.650 103.590 ;
        RECT 70.490 102.590 72.050 102.820 ;
        RECT 70.130 102.080 70.440 102.430 ;
        RECT 68.160 100.590 68.500 101.910 ;
        RECT 70.210 101.230 70.440 102.080 ;
        RECT 71.160 101.160 71.410 102.590 ;
        RECT 75.240 102.430 75.420 103.460 ;
        RECT 83.370 103.440 83.650 103.460 ;
        RECT 72.100 102.090 72.330 102.430 ;
        RECT 72.620 102.090 72.920 102.110 ;
        RECT 73.240 102.090 73.470 102.430 ;
        RECT 72.100 101.710 73.470 102.090 ;
        RECT 72.100 101.230 72.370 101.710 ;
        RECT 71.160 101.070 71.420 101.160 ;
        RECT 70.490 100.840 72.050 101.070 ;
        RECT 71.200 100.590 71.420 100.840 ;
        RECT 68.160 100.370 71.440 100.590 ;
        RECT 68.210 100.340 71.440 100.370 ;
        RECT 39.110 98.610 42.190 100.100 ;
        RECT 72.210 99.370 72.370 101.230 ;
        RECT 73.210 101.230 73.470 101.710 ;
        RECT 75.130 101.590 75.420 102.430 ;
        RECT 75.130 101.230 75.360 101.590 ;
        RECT 71.900 99.280 72.410 99.370 ;
        RECT 73.210 99.280 73.370 101.230 ;
        RECT 70.090 99.020 72.410 99.280 ;
        RECT 70.090 99.010 72.370 99.020 ;
        RECT 62.530 98.720 63.530 98.770 ;
        RECT 39.110 98.590 59.460 98.610 ;
        RECT 62.500 98.590 63.570 98.720 ;
        RECT 39.110 98.290 63.570 98.590 ;
        RECT 39.110 98.270 64.290 98.290 ;
        RECT 66.960 98.270 68.530 98.280 ;
        RECT 39.110 98.260 65.480 98.270 ;
        RECT 65.850 98.260 69.300 98.270 ;
        RECT 39.110 98.100 69.300 98.260 ;
        RECT 38.920 97.950 59.460 98.100 ;
        RECT 62.500 98.010 69.300 98.100 ;
        RECT 62.500 98.000 64.290 98.010 ;
        RECT 38.920 97.810 42.190 97.950 ;
        RECT 62.500 97.840 63.570 98.000 ;
        RECT 64.990 97.910 69.300 98.010 ;
        RECT 64.990 97.890 66.600 97.910 ;
        RECT 38.920 51.070 41.190 97.810 ;
        RECT 62.530 97.770 63.530 97.840 ;
        RECT 64.990 96.900 65.190 97.890 ;
        RECT 65.880 97.290 66.240 97.890 ;
        RECT 68.930 97.290 69.290 97.910 ;
        RECT 65.340 97.060 66.900 97.290 ;
        RECT 68.370 97.060 69.930 97.290 ;
        RECT 64.990 96.630 65.290 96.900 ;
        RECT 65.060 96.480 65.290 96.630 ;
        RECT 65.880 96.320 66.240 97.060 ;
        RECT 68.930 96.560 69.290 97.060 ;
        RECT 70.120 96.900 70.500 99.010 ;
        RECT 73.130 98.940 73.530 99.280 ;
        RECT 88.780 97.380 89.550 106.460 ;
        RECT 69.980 96.580 70.500 96.900 ;
        RECT 68.930 96.320 69.310 96.560 ;
        RECT 69.980 96.480 70.210 96.580 ;
        RECT 65.340 96.090 66.900 96.320 ;
        RECT 68.370 96.090 69.930 96.320 ;
        RECT 65.920 96.070 66.210 96.090 ;
        RECT 69.020 96.070 69.310 96.090 ;
        RECT 88.660 96.040 89.550 97.380 ;
        RECT 91.310 104.810 92.460 104.880 ;
        RECT 94.080 104.810 95.080 105.300 ;
        RECT 91.310 104.450 95.080 104.810 ;
        RECT 59.090 92.670 60.080 92.700 ;
        RECT 79.050 92.670 80.280 93.050 ;
        RECT 59.090 91.780 80.280 92.670 ;
        RECT 59.090 70.110 60.080 91.780 ;
        RECT 79.050 91.710 80.280 91.780 ;
        RECT 88.660 87.010 89.430 96.040 ;
        RECT 88.600 86.260 89.430 87.010 ;
        RECT 71.570 84.770 75.430 84.810 ;
        RECT 71.570 84.530 79.250 84.770 ;
        RECT 67.760 84.230 68.360 84.530 ;
        RECT 67.910 83.440 68.150 84.230 ;
        RECT 64.250 83.210 65.810 83.440 ;
        RECT 67.280 83.210 68.840 83.440 ;
        RECT 63.970 83.000 64.200 83.005 ;
        RECT 63.750 82.505 64.200 83.000 ;
        RECT 63.750 81.410 64.070 82.505 ;
        RECT 64.910 82.450 65.110 83.210 ;
        RECT 67.910 83.120 68.150 83.210 ;
        RECT 64.910 82.300 65.120 82.450 ;
        RECT 67.930 82.370 68.130 83.120 ;
        RECT 68.890 83.000 69.120 83.005 ;
        RECT 68.890 82.505 69.240 83.000 ;
        RECT 67.900 82.300 68.130 82.370 ;
        RECT 64.250 82.070 65.810 82.300 ;
        RECT 67.280 82.070 68.840 82.300 ;
        RECT 64.920 81.410 65.120 82.070 ;
        RECT 63.750 81.370 65.120 81.410 ;
        RECT 67.900 81.370 68.100 82.070 ;
        RECT 63.750 81.140 68.100 81.370 ;
        RECT 63.750 81.120 68.080 81.140 ;
        RECT 63.750 79.920 64.070 81.120 ;
        RECT 64.920 81.110 68.080 81.120 ;
        RECT 69.010 80.990 69.240 82.505 ;
        RECT 68.990 80.770 70.700 80.990 ;
        RECT 70.420 80.490 70.700 80.770 ;
        RECT 63.740 76.180 64.080 79.920 ;
        RECT 70.440 78.530 70.670 80.490 ;
        RECT 71.570 79.360 71.850 84.530 ;
        RECT 75.350 84.510 79.250 84.530 ;
        RECT 78.990 83.640 79.210 84.510 ;
        RECT 74.350 83.090 75.060 83.620 ;
        RECT 78.300 83.410 79.860 83.640 ;
        RECT 81.330 83.410 82.890 83.640 ;
        RECT 78.990 83.260 79.210 83.410 ;
        RECT 77.850 83.205 78.140 83.250 ;
        RECT 71.580 78.950 71.820 79.360 ;
        RECT 71.570 78.750 71.830 78.950 ;
        RECT 74.500 78.750 74.780 83.090 ;
        RECT 77.850 82.705 78.250 83.205 ;
        RECT 77.850 81.520 78.140 82.705 ;
        RECT 79.000 82.540 79.200 83.260 ;
        RECT 78.980 82.500 79.240 82.540 ;
        RECT 82.000 82.500 82.200 83.410 ;
        RECT 82.940 83.130 83.170 83.205 ;
        RECT 82.940 82.705 83.340 83.130 ;
        RECT 78.300 82.270 79.860 82.500 ;
        RECT 81.330 82.270 82.890 82.500 ;
        RECT 78.980 81.910 79.240 82.270 ;
        RECT 82.040 81.910 82.180 82.270 ;
        RECT 78.980 81.850 82.200 81.910 ;
        RECT 83.070 81.850 83.340 82.705 ;
        RECT 78.980 81.620 83.340 81.850 ;
        RECT 82.190 81.560 83.340 81.620 ;
        RECT 77.850 81.350 78.120 81.520 ;
        RECT 75.580 81.070 78.120 81.350 ;
        RECT 75.580 79.200 75.900 81.070 ;
        RECT 83.070 80.570 83.340 81.560 ;
        RECT 83.070 80.050 83.360 80.570 ;
        RECT 70.450 78.315 70.660 78.530 ;
        RECT 70.810 78.520 72.370 78.750 ;
        RECT 73.840 78.520 75.400 78.750 ;
        RECT 70.450 77.860 70.760 78.315 ;
        RECT 70.530 77.715 70.760 77.860 ;
        RECT 71.570 77.510 71.830 78.520 ;
        RECT 72.420 78.130 72.650 78.315 ;
        RECT 73.560 78.130 73.790 78.315 ;
        RECT 72.420 77.950 73.790 78.130 ;
        RECT 72.420 77.715 72.650 77.950 ;
        RECT 70.810 77.280 72.370 77.510 ;
        RECT 72.940 76.520 73.210 77.950 ;
        RECT 73.560 77.715 73.790 77.950 ;
        RECT 74.490 77.510 74.810 78.520 ;
        RECT 75.590 78.315 75.900 79.200 ;
        RECT 75.450 77.800 75.900 78.315 ;
        RECT 75.450 77.715 75.680 77.800 ;
        RECT 83.090 77.640 83.360 80.050 ;
        RECT 73.840 77.280 75.400 77.510 ;
        RECT 63.760 75.840 64.080 76.180 ;
        RECT 63.760 75.700 70.020 75.840 ;
        RECT 63.760 75.630 70.030 75.700 ;
        RECT 63.760 75.620 64.080 75.630 ;
        RECT 61.190 74.330 62.060 74.510 ;
        RECT 67.610 74.330 68.610 74.530 ;
        RECT 61.190 73.680 68.610 74.330 ;
        RECT 69.850 74.050 70.030 75.630 ;
        RECT 72.640 75.520 73.640 76.520 ;
        RECT 83.090 75.360 83.370 77.640 ;
        RECT 74.970 75.210 83.370 75.360 ;
        RECT 74.960 75.080 83.370 75.210 ;
        RECT 70.210 74.210 71.770 74.440 ;
        RECT 69.850 73.700 70.160 74.050 ;
        RECT 61.190 73.620 62.060 73.680 ;
        RECT 67.610 73.530 68.610 73.680 ;
        RECT 67.880 72.210 68.220 73.530 ;
        RECT 69.930 72.850 70.160 73.700 ;
        RECT 70.880 72.780 71.130 74.210 ;
        RECT 74.960 74.050 75.140 75.080 ;
        RECT 83.090 75.060 83.370 75.080 ;
        RECT 88.600 76.850 89.370 86.260 ;
        RECT 71.820 73.710 72.050 74.050 ;
        RECT 72.340 73.710 72.640 73.730 ;
        RECT 72.960 73.710 73.190 74.050 ;
        RECT 71.820 73.330 73.190 73.710 ;
        RECT 71.820 72.850 72.090 73.330 ;
        RECT 70.880 72.690 71.140 72.780 ;
        RECT 70.210 72.460 71.770 72.690 ;
        RECT 70.920 72.210 71.140 72.460 ;
        RECT 67.880 71.990 71.160 72.210 ;
        RECT 67.930 71.960 71.160 71.990 ;
        RECT 71.930 70.990 72.090 72.850 ;
        RECT 72.930 72.850 73.190 73.330 ;
        RECT 74.850 73.210 75.140 74.050 ;
        RECT 74.850 72.850 75.080 73.210 ;
        RECT 71.620 70.900 72.130 70.990 ;
        RECT 72.930 70.900 73.090 72.850 ;
        RECT 69.810 70.640 72.130 70.900 ;
        RECT 69.810 70.630 72.090 70.640 ;
        RECT 62.250 70.110 63.250 70.390 ;
        RECT 59.020 69.910 63.250 70.110 ;
        RECT 59.020 69.890 64.010 69.910 ;
        RECT 66.680 69.890 68.250 69.900 ;
        RECT 59.020 69.880 65.200 69.890 ;
        RECT 65.570 69.880 69.020 69.890 ;
        RECT 59.020 69.800 69.020 69.880 ;
        RECT 62.250 69.630 69.020 69.800 ;
        RECT 62.250 69.620 64.010 69.630 ;
        RECT 62.250 69.390 63.250 69.620 ;
        RECT 64.710 69.530 69.020 69.630 ;
        RECT 64.710 69.510 66.320 69.530 ;
        RECT 64.710 68.520 64.910 69.510 ;
        RECT 65.600 68.910 65.960 69.510 ;
        RECT 68.650 68.910 69.010 69.530 ;
        RECT 65.060 68.680 66.620 68.910 ;
        RECT 68.090 68.680 69.650 68.910 ;
        RECT 64.710 68.250 65.010 68.520 ;
        RECT 64.780 68.100 65.010 68.250 ;
        RECT 65.600 67.940 65.960 68.680 ;
        RECT 68.650 68.180 69.010 68.680 ;
        RECT 69.840 68.520 70.220 70.630 ;
        RECT 72.850 70.560 73.250 70.900 ;
        RECT 88.600 70.180 89.440 76.850 ;
        RECT 91.310 75.500 92.460 104.450 ;
        RECT 94.080 104.250 95.080 104.450 ;
        RECT 95.630 103.320 96.190 106.460 ;
        RECT 96.740 104.800 97.080 108.540 ;
        RECT 103.440 107.150 103.670 109.110 ;
        RECT 104.570 107.980 104.850 113.150 ;
        RECT 108.350 113.130 112.250 113.150 ;
        RECT 111.990 112.260 112.210 113.130 ;
        RECT 107.350 111.710 108.060 112.240 ;
        RECT 111.300 112.030 112.860 112.260 ;
        RECT 114.330 112.030 115.890 112.260 ;
        RECT 111.990 111.880 112.210 112.030 ;
        RECT 110.850 111.825 111.140 111.870 ;
        RECT 104.580 107.570 104.820 107.980 ;
        RECT 104.570 107.370 104.830 107.570 ;
        RECT 107.500 107.370 107.780 111.710 ;
        RECT 110.850 111.325 111.250 111.825 ;
        RECT 110.850 110.140 111.140 111.325 ;
        RECT 112.000 111.160 112.200 111.880 ;
        RECT 111.980 111.120 112.240 111.160 ;
        RECT 115.000 111.120 115.200 112.030 ;
        RECT 115.940 111.750 116.170 111.825 ;
        RECT 115.940 111.325 116.340 111.750 ;
        RECT 111.300 110.890 112.860 111.120 ;
        RECT 114.330 110.890 115.890 111.120 ;
        RECT 111.980 110.530 112.240 110.890 ;
        RECT 115.040 110.530 115.180 110.890 ;
        RECT 111.980 110.470 115.200 110.530 ;
        RECT 116.070 110.470 116.340 111.325 ;
        RECT 111.980 110.240 116.340 110.470 ;
        RECT 115.190 110.180 116.340 110.240 ;
        RECT 110.850 109.970 111.120 110.140 ;
        RECT 108.580 109.690 111.120 109.970 ;
        RECT 108.580 107.820 108.900 109.690 ;
        RECT 116.070 109.190 116.340 110.180 ;
        RECT 116.070 108.670 116.360 109.190 ;
        RECT 103.450 106.935 103.660 107.150 ;
        RECT 103.810 107.140 105.370 107.370 ;
        RECT 106.840 107.140 108.400 107.370 ;
        RECT 103.450 106.480 103.760 106.935 ;
        RECT 103.530 106.335 103.760 106.480 ;
        RECT 104.570 106.130 104.830 107.140 ;
        RECT 105.420 106.750 105.650 106.935 ;
        RECT 106.560 106.750 106.790 106.935 ;
        RECT 105.420 106.570 106.790 106.750 ;
        RECT 105.420 106.335 105.650 106.570 ;
        RECT 103.810 105.900 105.370 106.130 ;
        RECT 105.940 105.140 106.210 106.570 ;
        RECT 106.560 106.335 106.790 106.570 ;
        RECT 107.490 106.130 107.810 107.140 ;
        RECT 108.590 106.935 108.900 107.820 ;
        RECT 108.450 106.420 108.900 106.935 ;
        RECT 108.450 106.335 108.680 106.420 ;
        RECT 116.090 106.260 116.360 108.670 ;
        RECT 106.840 105.900 108.400 106.130 ;
        RECT 96.760 104.460 97.080 104.800 ;
        RECT 96.760 104.320 103.020 104.460 ;
        RECT 96.760 104.250 103.030 104.320 ;
        RECT 96.760 104.240 97.080 104.250 ;
        RECT 95.790 102.960 96.190 103.320 ;
        RECT 100.610 102.960 101.610 103.150 ;
        RECT 95.790 102.270 101.610 102.960 ;
        RECT 102.850 102.670 103.030 104.250 ;
        RECT 105.640 104.140 106.640 105.140 ;
        RECT 116.090 103.980 116.370 106.260 ;
        RECT 107.970 103.830 116.370 103.980 ;
        RECT 107.960 103.700 116.370 103.830 ;
        RECT 103.210 102.830 104.770 103.060 ;
        RECT 106.240 102.830 107.800 103.060 ;
        RECT 102.850 102.320 103.160 102.670 ;
        RECT 100.610 102.150 101.610 102.270 ;
        RECT 100.880 100.830 101.220 102.150 ;
        RECT 102.930 101.470 103.160 102.320 ;
        RECT 103.880 101.400 104.130 102.830 ;
        RECT 104.820 102.330 105.050 102.670 ;
        RECT 105.340 102.330 105.640 102.350 ;
        RECT 105.960 102.330 106.190 102.670 ;
        RECT 104.820 101.950 106.190 102.330 ;
        RECT 104.820 101.470 105.090 101.950 ;
        RECT 103.880 101.310 104.140 101.400 ;
        RECT 103.210 101.080 104.770 101.310 ;
        RECT 103.920 100.830 104.140 101.080 ;
        RECT 100.880 100.610 104.160 100.830 ;
        RECT 100.930 100.580 104.160 100.610 ;
        RECT 104.930 99.610 105.090 101.470 ;
        RECT 105.930 101.470 106.190 101.950 ;
        RECT 106.860 101.470 107.110 102.830 ;
        RECT 107.960 102.670 108.140 103.700 ;
        RECT 116.090 103.680 116.370 103.700 ;
        RECT 136.640 104.940 139.250 137.860 ;
        RECT 107.850 101.830 108.140 102.670 ;
        RECT 109.760 101.980 110.760 102.980 ;
        RECT 107.850 101.470 108.080 101.830 ;
        RECT 104.620 99.520 105.130 99.610 ;
        RECT 105.930 99.520 106.090 101.470 ;
        RECT 106.860 101.310 107.120 101.470 ;
        RECT 106.240 101.080 107.800 101.310 ;
        RECT 110.080 101.250 110.450 101.980 ;
        RECT 106.890 100.560 107.120 101.080 ;
        RECT 110.080 100.750 110.460 101.250 ;
        RECT 136.640 100.750 138.930 104.940 ;
        RECT 109.820 100.560 138.930 100.750 ;
        RECT 106.890 100.270 138.930 100.560 ;
        RECT 109.820 100.260 138.930 100.270 ;
        RECT 110.080 100.230 110.460 100.260 ;
        RECT 136.640 100.030 138.930 100.260 ;
        RECT 102.810 99.260 105.130 99.520 ;
        RECT 102.810 99.250 105.090 99.260 ;
        RECT 95.250 98.530 96.250 99.010 ;
        RECT 95.250 98.510 97.010 98.530 ;
        RECT 99.680 98.510 101.250 98.520 ;
        RECT 95.250 98.500 98.200 98.510 ;
        RECT 98.570 98.500 102.020 98.510 ;
        RECT 95.250 98.250 102.020 98.500 ;
        RECT 95.250 98.240 97.010 98.250 ;
        RECT 95.250 98.010 96.250 98.240 ;
        RECT 97.710 98.150 102.020 98.250 ;
        RECT 97.710 98.130 99.320 98.150 ;
        RECT 97.710 97.140 97.910 98.130 ;
        RECT 98.600 97.530 98.960 98.130 ;
        RECT 101.650 97.530 102.010 98.150 ;
        RECT 98.060 97.300 99.620 97.530 ;
        RECT 101.090 97.300 102.650 97.530 ;
        RECT 97.710 96.870 98.010 97.140 ;
        RECT 97.780 96.720 98.010 96.870 ;
        RECT 98.600 96.560 98.960 97.300 ;
        RECT 101.650 96.800 102.010 97.300 ;
        RECT 102.840 97.140 103.220 99.250 ;
        RECT 105.850 99.180 106.250 99.520 ;
        RECT 102.700 96.820 103.220 97.140 ;
        RECT 101.650 96.560 102.030 96.800 ;
        RECT 102.700 96.720 102.930 96.820 ;
        RECT 98.060 96.330 99.620 96.560 ;
        RECT 101.090 96.330 102.650 96.560 ;
        RECT 98.640 96.310 98.930 96.330 ;
        RECT 101.740 96.310 102.030 96.330 ;
        RECT 103.220 87.290 107.080 87.330 ;
        RECT 103.220 87.050 110.900 87.290 ;
        RECT 99.410 86.750 100.010 87.050 ;
        RECT 99.560 85.960 99.800 86.750 ;
        RECT 95.900 85.730 97.460 85.960 ;
        RECT 98.930 85.730 100.490 85.960 ;
        RECT 95.620 85.520 95.850 85.525 ;
        RECT 95.400 85.025 95.850 85.520 ;
        RECT 95.400 83.930 95.720 85.025 ;
        RECT 96.560 84.970 96.760 85.730 ;
        RECT 99.560 85.640 99.800 85.730 ;
        RECT 96.560 84.820 96.770 84.970 ;
        RECT 99.580 84.890 99.780 85.640 ;
        RECT 100.540 85.520 100.770 85.525 ;
        RECT 100.540 85.025 100.890 85.520 ;
        RECT 99.550 84.820 99.780 84.890 ;
        RECT 95.900 84.590 97.460 84.820 ;
        RECT 98.930 84.590 100.490 84.820 ;
        RECT 96.570 83.930 96.770 84.590 ;
        RECT 95.400 83.890 96.770 83.930 ;
        RECT 99.550 83.890 99.750 84.590 ;
        RECT 95.400 83.660 99.750 83.890 ;
        RECT 95.400 83.640 99.730 83.660 ;
        RECT 95.400 82.440 95.720 83.640 ;
        RECT 96.570 83.630 99.730 83.640 ;
        RECT 100.660 83.510 100.890 85.025 ;
        RECT 100.640 83.290 102.350 83.510 ;
        RECT 102.070 83.010 102.350 83.290 ;
        RECT 95.390 78.700 95.730 82.440 ;
        RECT 102.090 81.050 102.320 83.010 ;
        RECT 103.220 81.880 103.500 87.050 ;
        RECT 107.000 87.030 110.900 87.050 ;
        RECT 110.640 86.160 110.860 87.030 ;
        RECT 106.000 85.610 106.710 86.140 ;
        RECT 109.950 85.930 111.510 86.160 ;
        RECT 112.980 85.930 114.540 86.160 ;
        RECT 110.640 85.780 110.860 85.930 ;
        RECT 109.500 85.725 109.790 85.770 ;
        RECT 103.230 81.470 103.470 81.880 ;
        RECT 103.220 81.270 103.480 81.470 ;
        RECT 106.150 81.270 106.430 85.610 ;
        RECT 109.500 85.225 109.900 85.725 ;
        RECT 109.500 84.040 109.790 85.225 ;
        RECT 110.650 85.060 110.850 85.780 ;
        RECT 110.630 85.020 110.890 85.060 ;
        RECT 113.650 85.020 113.850 85.930 ;
        RECT 114.590 85.650 114.820 85.725 ;
        RECT 114.590 85.225 114.990 85.650 ;
        RECT 109.950 84.790 111.510 85.020 ;
        RECT 112.980 84.790 114.540 85.020 ;
        RECT 110.630 84.430 110.890 84.790 ;
        RECT 113.690 84.430 113.830 84.790 ;
        RECT 110.630 84.370 113.850 84.430 ;
        RECT 114.720 84.370 114.990 85.225 ;
        RECT 110.630 84.140 114.990 84.370 ;
        RECT 113.840 84.080 114.990 84.140 ;
        RECT 109.500 83.870 109.770 84.040 ;
        RECT 107.230 83.590 109.770 83.870 ;
        RECT 107.230 81.720 107.550 83.590 ;
        RECT 114.720 83.090 114.990 84.080 ;
        RECT 114.720 82.570 115.010 83.090 ;
        RECT 102.100 80.835 102.310 81.050 ;
        RECT 102.460 81.040 104.020 81.270 ;
        RECT 105.490 81.040 107.050 81.270 ;
        RECT 102.100 80.380 102.410 80.835 ;
        RECT 102.180 80.235 102.410 80.380 ;
        RECT 103.220 80.030 103.480 81.040 ;
        RECT 104.070 80.650 104.300 80.835 ;
        RECT 105.210 80.650 105.440 80.835 ;
        RECT 104.070 80.470 105.440 80.650 ;
        RECT 104.070 80.235 104.300 80.470 ;
        RECT 102.460 79.800 104.020 80.030 ;
        RECT 104.590 79.040 104.860 80.470 ;
        RECT 105.210 80.235 105.440 80.470 ;
        RECT 106.140 80.030 106.460 81.040 ;
        RECT 107.240 80.835 107.550 81.720 ;
        RECT 107.100 80.320 107.550 80.835 ;
        RECT 107.100 80.235 107.330 80.320 ;
        RECT 114.740 80.160 115.010 82.570 ;
        RECT 105.490 79.800 107.050 80.030 ;
        RECT 95.410 78.360 95.730 78.700 ;
        RECT 95.410 78.220 101.670 78.360 ;
        RECT 95.410 78.150 101.680 78.220 ;
        RECT 95.410 78.140 95.730 78.150 ;
        RECT 99.260 76.850 100.260 77.050 ;
        RECT 99.230 76.060 100.260 76.850 ;
        RECT 101.500 76.570 101.680 78.150 ;
        RECT 104.290 78.040 105.290 79.040 ;
        RECT 114.740 77.880 115.020 80.160 ;
        RECT 106.620 77.730 115.020 77.880 ;
        RECT 106.610 77.600 115.020 77.730 ;
        RECT 101.860 76.730 103.420 76.960 ;
        RECT 104.890 76.730 106.450 76.960 ;
        RECT 101.500 76.220 101.810 76.570 ;
        RECT 99.260 76.050 100.260 76.060 ;
        RECT 91.480 72.810 92.460 75.500 ;
        RECT 99.530 74.730 99.870 76.050 ;
        RECT 101.580 75.370 101.810 76.220 ;
        RECT 102.530 75.300 102.780 76.730 ;
        RECT 103.470 76.230 103.700 76.570 ;
        RECT 103.990 76.230 104.290 76.250 ;
        RECT 104.610 76.230 104.840 76.570 ;
        RECT 103.470 75.850 104.840 76.230 ;
        RECT 103.470 75.370 103.740 75.850 ;
        RECT 102.530 75.210 102.790 75.300 ;
        RECT 101.860 74.980 103.420 75.210 ;
        RECT 102.570 74.730 102.790 74.980 ;
        RECT 99.530 74.510 102.810 74.730 ;
        RECT 99.580 74.480 102.810 74.510 ;
        RECT 103.580 73.510 103.740 75.370 ;
        RECT 104.580 75.370 104.840 75.850 ;
        RECT 105.510 75.370 105.760 76.730 ;
        RECT 106.610 76.570 106.790 77.600 ;
        RECT 114.740 77.580 115.020 77.600 ;
        RECT 106.500 75.730 106.790 76.570 ;
        RECT 108.410 76.810 109.410 76.880 ;
        RECT 136.730 76.810 138.820 100.030 ;
        RECT 108.410 75.880 138.930 76.810 ;
        RECT 106.500 75.370 106.730 75.730 ;
        RECT 103.270 73.420 103.780 73.510 ;
        RECT 104.580 73.420 104.740 75.370 ;
        RECT 105.510 75.210 105.770 75.370 ;
        RECT 104.890 74.980 106.450 75.210 ;
        RECT 108.730 75.150 109.100 75.880 ;
        RECT 105.540 74.460 105.770 74.980 ;
        RECT 108.730 74.460 109.110 75.150 ;
        RECT 105.540 74.170 109.110 74.460 ;
        RECT 108.730 74.130 109.110 74.170 ;
        RECT 101.460 73.160 103.780 73.420 ;
        RECT 101.460 73.150 103.740 73.160 ;
        RECT 93.900 72.810 94.900 72.910 ;
        RECT 91.480 72.430 95.220 72.810 ;
        RECT 91.480 72.410 95.660 72.430 ;
        RECT 98.330 72.410 99.900 72.420 ;
        RECT 91.480 72.400 96.850 72.410 ;
        RECT 97.220 72.400 100.670 72.410 ;
        RECT 91.480 72.160 100.670 72.400 ;
        RECT 91.480 72.060 92.460 72.160 ;
        RECT 93.900 72.150 100.670 72.160 ;
        RECT 93.900 72.140 95.660 72.150 ;
        RECT 93.900 71.910 94.900 72.140 ;
        RECT 96.360 72.050 100.670 72.150 ;
        RECT 96.360 72.030 97.970 72.050 ;
        RECT 96.360 71.040 96.560 72.030 ;
        RECT 97.250 71.430 97.610 72.030 ;
        RECT 100.300 71.430 100.660 72.050 ;
        RECT 96.710 71.200 98.270 71.430 ;
        RECT 99.740 71.200 101.300 71.430 ;
        RECT 96.360 70.770 96.660 71.040 ;
        RECT 96.430 70.620 96.660 70.770 ;
        RECT 97.250 70.460 97.610 71.200 ;
        RECT 100.300 70.700 100.660 71.200 ;
        RECT 101.490 71.040 101.870 73.150 ;
        RECT 104.500 73.080 104.900 73.420 ;
        RECT 101.350 70.720 101.870 71.040 ;
        RECT 100.300 70.460 100.680 70.700 ;
        RECT 101.350 70.620 101.580 70.720 ;
        RECT 96.710 70.230 98.270 70.460 ;
        RECT 99.740 70.230 101.300 70.460 ;
        RECT 97.290 70.210 97.580 70.230 ;
        RECT 100.390 70.210 100.680 70.230 ;
        RECT 88.600 69.050 93.730 70.180 ;
        RECT 69.700 68.200 70.220 68.520 ;
        RECT 68.650 67.940 69.030 68.180 ;
        RECT 69.700 68.100 69.930 68.200 ;
        RECT 65.060 67.710 66.620 67.940 ;
        RECT 68.090 67.710 69.650 67.940 ;
        RECT 65.640 67.690 65.930 67.710 ;
        RECT 68.740 67.690 69.030 67.710 ;
        RECT 91.430 63.550 92.050 63.780 ;
        RECT 85.380 63.100 86.970 63.340 ;
        RECT 73.100 62.410 86.970 63.100 ;
        RECT 73.110 61.100 73.760 62.410 ;
        RECT 85.380 61.940 86.970 62.410 ;
        RECT 90.980 62.400 92.470 63.550 ;
        RECT 91.430 61.830 92.050 62.400 ;
        RECT 87.590 61.370 92.050 61.830 ;
        RECT 72.910 60.100 73.910 61.100 ;
        RECT 75.180 61.020 76.180 61.370 ;
        RECT 87.560 61.070 92.050 61.370 ;
        RECT 75.180 60.590 78.870 61.020 ;
        RECT 75.180 60.370 76.180 60.590 ;
        RECT 73.180 59.170 73.490 60.100 ;
        RECT 72.590 58.940 74.150 59.170 ;
        RECT 73.110 58.930 73.490 58.940 ;
        RECT 72.310 58.720 72.540 58.780 ;
        RECT 73.110 58.750 73.420 58.930 ;
        RECT 75.240 58.780 75.480 60.370 ;
        RECT 75.620 58.940 77.180 59.170 ;
        RECT 72.020 58.280 72.540 58.720 ;
        RECT 73.020 58.660 73.540 58.750 ;
        RECT 74.200 58.660 74.430 58.780 ;
        RECT 73.020 58.440 74.430 58.660 ;
        RECT 73.020 58.330 73.540 58.440 ;
        RECT 72.020 56.710 72.400 58.280 ;
        RECT 73.110 58.120 73.420 58.330 ;
        RECT 74.200 58.280 74.430 58.440 ;
        RECT 75.240 58.430 75.570 58.780 ;
        RECT 76.240 58.750 76.550 58.940 ;
        RECT 75.340 58.280 75.570 58.430 ;
        RECT 76.100 58.330 76.620 58.750 ;
        RECT 77.230 58.630 77.460 58.780 ;
        RECT 76.240 58.120 76.550 58.330 ;
        RECT 77.230 58.280 77.670 58.630 ;
        RECT 72.590 57.890 74.150 58.120 ;
        RECT 75.620 57.890 77.180 58.120 ;
        RECT 72.590 56.870 74.150 57.100 ;
        RECT 75.620 56.870 77.180 57.100 ;
        RECT 72.020 56.590 72.540 56.710 ;
        RECT 73.160 56.610 73.500 56.870 ;
        RECT 76.170 56.670 76.480 56.870 ;
        RECT 77.360 56.710 77.670 58.280 ;
        RECT 72.900 56.600 73.500 56.610 ;
        RECT 72.860 56.590 73.550 56.600 ;
        RECT 72.020 56.310 73.550 56.590 ;
        RECT 72.020 56.230 72.540 56.310 ;
        RECT 72.860 56.300 73.550 56.310 ;
        RECT 72.310 56.210 72.540 56.230 ;
        RECT 73.160 56.050 73.500 56.300 ;
        RECT 76.110 56.290 76.610 56.670 ;
        RECT 76.170 56.050 76.480 56.290 ;
        RECT 77.230 56.270 77.670 56.710 ;
        RECT 77.230 56.210 77.460 56.270 ;
        RECT 72.590 55.820 74.150 56.050 ;
        RECT 75.620 55.820 77.180 56.050 ;
        RECT 78.280 53.090 78.840 60.590 ;
        RECT 87.560 59.940 88.220 61.070 ;
        RECT 91.430 61.010 92.050 61.070 ;
        RECT 89.590 60.050 90.590 60.210 ;
        RECT 87.320 58.940 88.320 59.940 ;
        RECT 89.590 59.290 93.640 60.050 ;
        RECT 89.590 59.210 90.590 59.290 ;
        RECT 87.590 58.010 87.900 58.940 ;
        RECT 87.000 57.780 88.560 58.010 ;
        RECT 87.520 57.770 87.900 57.780 ;
        RECT 86.720 57.560 86.950 57.620 ;
        RECT 87.520 57.590 87.830 57.770 ;
        RECT 89.650 57.620 89.890 59.210 ;
        RECT 90.030 57.780 91.590 58.010 ;
        RECT 86.430 57.120 86.950 57.560 ;
        RECT 87.430 57.500 87.950 57.590 ;
        RECT 88.610 57.500 88.840 57.620 ;
        RECT 87.430 57.280 88.840 57.500 ;
        RECT 87.430 57.170 87.950 57.280 ;
        RECT 86.430 55.550 86.810 57.120 ;
        RECT 87.520 56.960 87.830 57.170 ;
        RECT 88.610 57.120 88.840 57.280 ;
        RECT 89.650 57.270 89.980 57.620 ;
        RECT 90.650 57.590 90.960 57.780 ;
        RECT 89.750 57.120 89.980 57.270 ;
        RECT 90.510 57.170 91.030 57.590 ;
        RECT 91.640 57.470 91.870 57.620 ;
        RECT 90.650 56.960 90.960 57.170 ;
        RECT 91.640 57.120 92.080 57.470 ;
        RECT 87.000 56.730 88.560 56.960 ;
        RECT 90.030 56.730 91.590 56.960 ;
        RECT 87.000 55.710 88.560 55.940 ;
        RECT 90.030 55.710 91.590 55.940 ;
        RECT 86.430 55.430 86.950 55.550 ;
        RECT 87.570 55.450 87.910 55.710 ;
        RECT 90.580 55.510 90.890 55.710 ;
        RECT 91.770 55.550 92.080 57.120 ;
        RECT 87.310 55.440 87.910 55.450 ;
        RECT 87.270 55.430 87.960 55.440 ;
        RECT 86.430 55.150 87.960 55.430 ;
        RECT 86.430 55.070 86.950 55.150 ;
        RECT 87.270 55.140 87.960 55.150 ;
        RECT 86.720 55.050 86.950 55.070 ;
        RECT 87.570 54.890 87.910 55.140 ;
        RECT 90.520 55.130 91.020 55.510 ;
        RECT 90.580 54.890 90.890 55.130 ;
        RECT 91.640 55.110 92.080 55.550 ;
        RECT 91.640 55.050 91.870 55.110 ;
        RECT 87.000 54.660 88.560 54.890 ;
        RECT 90.030 54.660 91.590 54.890 ;
        RECT 78.280 52.720 78.900 53.090 ;
        RECT 38.920 50.380 41.130 51.070 ;
        RECT 38.790 49.550 41.130 50.380 ;
        RECT 38.600 47.090 41.130 49.550 ;
        RECT 78.340 41.950 78.900 52.720 ;
        RECT 82.560 47.330 83.860 47.590 ;
        RECT 81.290 46.550 84.730 47.330 ;
        RECT 81.320 43.370 81.640 46.550 ;
        RECT 82.560 46.460 83.860 46.550 ;
        RECT 84.370 43.370 84.690 46.550 ;
        RECT 80.770 43.140 82.330 43.370 ;
        RECT 83.800 43.140 85.360 43.370 ;
        RECT 81.320 43.080 81.640 43.140 ;
        RECT 80.490 42.770 80.720 42.935 ;
        RECT 80.030 42.570 80.720 42.770 ;
        RECT 78.130 41.710 79.130 41.950 ;
        RECT 80.030 41.710 80.190 42.570 ;
        RECT 80.490 42.435 80.720 42.570 ;
        RECT 81.380 42.230 81.570 43.080 ;
        RECT 84.370 42.960 84.690 43.140 ;
        RECT 84.440 42.230 84.630 42.960 ;
        RECT 85.410 42.720 85.640 42.935 ;
        RECT 85.410 42.560 86.270 42.720 ;
        RECT 85.410 42.435 85.640 42.560 ;
        RECT 80.770 42.200 82.330 42.230 ;
        RECT 78.130 41.240 80.190 41.710 ;
        RECT 78.130 40.950 79.130 41.240 ;
        RECT 80.030 39.970 80.190 41.240 ;
        RECT 80.450 42.010 82.330 42.200 ;
        RECT 80.450 40.775 80.600 42.010 ;
        RECT 80.770 42.000 82.330 42.010 ;
        RECT 83.800 42.180 85.360 42.230 ;
        RECT 83.800 42.020 85.740 42.180 ;
        RECT 83.800 42.000 85.360 42.020 ;
        RECT 80.770 40.980 82.330 41.210 ;
        RECT 83.800 40.980 85.360 41.210 ;
        RECT 80.450 40.420 80.720 40.775 ;
        RECT 80.490 40.275 80.720 40.420 ;
        RECT 81.360 40.070 81.550 40.980 ;
        RECT 84.430 40.070 84.620 40.980 ;
        RECT 85.540 40.775 85.720 42.020 ;
        RECT 85.410 40.400 85.720 40.775 ;
        RECT 86.020 41.310 86.270 42.560 ;
        RECT 86.880 41.540 87.880 41.620 ;
        RECT 92.630 41.540 93.640 59.290 ;
        RECT 86.880 41.310 93.640 41.540 ;
        RECT 86.020 40.840 93.640 41.310 ;
        RECT 85.410 40.275 85.640 40.400 ;
        RECT 80.770 39.970 82.330 40.070 ;
        RECT 80.030 39.840 82.330 39.970 ;
        RECT 83.800 40.040 85.360 40.070 ;
        RECT 86.020 40.040 86.270 40.840 ;
        RECT 86.880 40.720 93.640 40.840 ;
        RECT 86.880 40.620 87.880 40.720 ;
        RECT 83.800 39.890 86.270 40.040 ;
        RECT 83.800 39.880 86.090 39.890 ;
        RECT 83.800 39.840 85.360 39.880 ;
        RECT 80.030 39.830 81.390 39.840 ;
      LAYER met2 ;
        RECT 101.420 212.190 101.740 212.270 ;
        RECT 101.400 211.730 101.740 212.190 ;
        RECT 94.530 210.020 95.110 210.670 ;
        RECT 98.310 210.070 98.730 210.660 ;
        RECT 99.340 209.960 99.950 210.690 ;
        RECT 101.400 210.620 101.700 211.730 ;
        RECT 101.400 210.080 101.720 210.620 ;
        RECT 101.450 209.540 101.610 210.080 ;
        RECT 103.160 210.010 103.770 210.740 ;
        RECT 101.430 209.490 101.690 209.540 ;
        RECT 96.540 209.130 101.690 209.490 ;
        RECT 74.280 208.850 74.590 208.920 ;
        RECT 78.530 208.850 78.890 208.930 ;
        RECT 96.540 208.920 96.740 209.130 ;
        RECT 101.430 209.090 101.690 209.130 ;
        RECT 74.170 208.630 78.890 208.850 ;
        RECT 74.280 208.480 74.590 208.630 ;
        RECT 78.530 208.550 78.890 208.630 ;
        RECT 96.550 208.530 96.700 208.920 ;
        RECT 96.520 208.050 96.780 208.530 ;
        RECT 94.520 206.360 95.010 206.950 ;
        RECT 96.600 206.930 96.760 208.050 ;
        RECT 101.410 208.000 101.680 208.490 ;
        RECT 96.530 206.450 96.790 206.930 ;
        RECT 98.320 206.370 98.810 206.960 ;
        RECT 99.460 206.430 99.950 207.020 ;
        RECT 101.480 206.910 101.620 208.000 ;
        RECT 101.430 206.420 101.700 206.910 ;
        RECT 101.460 205.850 101.650 206.420 ;
        RECT 103.220 206.390 103.710 206.980 ;
        RECT 101.350 205.810 101.670 205.850 ;
        RECT 96.510 205.520 101.670 205.810 ;
        RECT 96.510 205.390 96.740 205.520 ;
        RECT 101.350 205.450 101.670 205.520 ;
        RECT 96.540 204.910 96.740 205.390 ;
        RECT 96.480 204.300 96.780 204.910 ;
        RECT 94.490 202.680 95.000 203.340 ;
        RECT 96.530 203.310 96.720 204.300 ;
        RECT 96.490 202.700 96.790 203.310 ;
        RECT 98.320 202.680 98.830 203.340 ;
        RECT 99.430 202.670 99.920 203.370 ;
        RECT 103.230 202.700 103.720 203.400 ;
        RECT 143.400 187.080 143.760 187.110 ;
        RECT 121.190 186.460 143.760 187.080 ;
        RECT 121.190 186.220 121.890 186.460 ;
        RECT 121.110 185.130 121.890 186.220 ;
        RECT 131.300 185.920 131.760 185.980 ;
        RECT 121.190 185.000 121.890 185.130 ;
        RECT 131.090 185.900 131.870 185.920 ;
        RECT 131.090 185.690 131.880 185.900 ;
        RECT 131.090 185.200 131.990 185.690 ;
        RECT 131.090 185.100 131.880 185.200 ;
        RECT 110.930 184.260 111.520 184.370 ;
        RECT 91.240 183.980 91.780 184.080 ;
        RECT 86.000 183.400 91.810 183.980 ;
        RECT 105.700 183.760 111.640 184.260 ;
        RECT 46.170 181.610 46.580 181.690 ;
        RECT 56.810 181.620 57.390 181.880 ;
        RECT 55.710 181.610 57.390 181.620 ;
        RECT 46.070 181.460 57.390 181.610 ;
        RECT 46.170 181.340 57.390 181.460 ;
        RECT 46.170 181.330 47.960 181.340 ;
        RECT 46.170 181.190 46.580 181.330 ;
        RECT 47.660 180.400 47.960 181.330 ;
        RECT 55.710 181.290 57.390 181.340 ;
        RECT 56.810 181.060 57.390 181.290 ;
        RECT 67.720 181.380 68.100 181.520 ;
        RECT 68.930 181.380 69.200 181.530 ;
        RECT 67.720 181.150 69.200 181.380 ;
        RECT 67.720 181.010 68.100 181.150 ;
        RECT 47.610 179.900 47.990 180.400 ;
        RECT 47.660 178.810 47.960 179.900 ;
        RECT 47.610 178.310 47.990 178.810 ;
        RECT 47.660 177.260 47.960 178.310 ;
        RECT 64.270 178.260 64.720 178.450 ;
        RECT 60.180 178.150 65.740 178.260 ;
        RECT 67.700 178.150 68.080 178.240 ;
        RECT 60.180 177.980 68.080 178.150 ;
        RECT 60.180 177.770 60.830 177.980 ;
        RECT 64.270 177.940 68.080 177.980 ;
        RECT 64.270 177.810 64.720 177.940 ;
        RECT 67.700 177.800 68.080 177.940 ;
        RECT 68.920 177.800 69.200 181.150 ;
        RECT 70.070 181.310 70.340 181.470 ;
        RECT 71.750 181.460 76.190 181.470 ;
        RECT 71.720 181.400 76.190 181.460 ;
        RECT 86.000 181.400 86.550 183.400 ;
        RECT 71.720 181.310 86.550 181.400 ;
        RECT 70.070 181.070 86.550 181.310 ;
        RECT 70.070 180.980 70.340 181.070 ;
        RECT 71.720 181.040 86.550 181.070 ;
        RECT 71.720 180.940 71.980 181.040 ;
        RECT 76.930 181.000 86.550 181.040 ;
        RECT 86.000 180.970 86.550 181.000 ;
        RECT 89.540 181.310 89.910 181.480 ;
        RECT 90.770 181.310 91.050 181.420 ;
        RECT 89.540 181.100 91.050 181.310 ;
        RECT 89.540 180.910 89.910 181.100 ;
        RECT 90.770 181.010 91.050 181.100 ;
        RECT 91.780 181.300 92.180 181.470 ;
        RECT 93.080 181.300 93.350 181.440 ;
        RECT 91.780 181.140 93.350 181.300 ;
        RECT 91.780 181.030 92.180 181.140 ;
        RECT 93.080 181.010 93.350 181.140 ;
        RECT 90.140 180.700 90.520 180.840 ;
        RECT 91.350 180.700 91.620 180.850 ;
        RECT 90.140 180.470 91.620 180.700 ;
        RECT 90.140 180.330 90.520 180.470 ;
        RECT 69.960 177.990 70.460 178.210 ;
        RECT 73.430 177.990 73.740 178.060 ;
        RECT 47.650 176.680 48.030 177.260 ;
        RECT 47.660 175.670 47.960 176.680 ;
        RECT 47.630 175.090 48.010 175.670 ;
        RECT 47.660 174.800 47.960 175.090 ;
        RECT 47.660 174.050 48.010 174.800 ;
        RECT 47.660 173.470 48.050 174.050 ;
        RECT 47.660 172.450 48.010 173.470 ;
        RECT 47.610 171.870 48.010 172.450 ;
        RECT 47.660 170.840 48.010 171.870 ;
        RECT 47.630 170.310 48.030 170.840 ;
        RECT 47.680 169.190 47.960 170.310 ;
        RECT 47.650 168.690 48.030 169.190 ;
        RECT 47.680 167.610 47.960 168.690 ;
        RECT 47.610 167.110 47.990 167.610 ;
        RECT 47.680 166.030 47.960 167.110 ;
        RECT 47.640 165.530 48.020 166.030 ;
        RECT 47.720 160.030 47.960 165.530 ;
        RECT 46.460 159.880 46.890 159.990 ;
        RECT 47.630 159.880 48.060 160.030 ;
        RECT 46.460 159.590 48.060 159.880 ;
        RECT 46.460 159.410 46.890 159.590 ;
        RECT 47.630 159.450 48.060 159.590 ;
        RECT 47.040 159.090 47.470 159.190 ;
        RECT 48.230 159.090 48.660 159.190 ;
        RECT 47.040 158.990 48.660 159.090 ;
        RECT 47.040 158.800 48.910 158.990 ;
        RECT 47.040 158.610 47.470 158.800 ;
        RECT 48.230 158.610 48.910 158.800 ;
        RECT 46.480 157.030 46.890 157.240 ;
        RECT 47.700 157.030 48.110 157.300 ;
        RECT 46.480 156.860 48.110 157.030 ;
        RECT 46.480 156.740 46.890 156.860 ;
        RECT 47.700 156.800 48.110 156.860 ;
        RECT 47.110 156.230 47.520 156.430 ;
        RECT 48.410 156.380 48.910 158.610 ;
        RECT 48.290 156.230 48.910 156.380 ;
        RECT 47.110 156.060 48.910 156.230 ;
        RECT 47.110 155.930 47.520 156.060 ;
        RECT 48.290 155.880 48.910 156.060 ;
        RECT 48.410 155.860 48.910 155.880 ;
        RECT 60.140 153.190 60.830 177.770 ;
        RECT 67.020 177.590 67.510 177.630 ;
        RECT 68.280 177.590 68.610 177.680 ;
        RECT 67.020 177.330 68.700 177.590 ;
        RECT 67.020 177.310 68.610 177.330 ;
        RECT 67.020 177.080 67.510 177.310 ;
        RECT 68.280 177.220 68.610 177.310 ;
        RECT 68.920 177.210 69.220 177.800 ;
        RECT 69.960 177.550 79.150 177.990 ;
        RECT 81.780 177.700 82.770 177.720 ;
        RECT 81.780 177.690 82.830 177.700 ;
        RECT 86.690 177.690 87.140 177.770 ;
        RECT 69.960 177.460 70.460 177.550 ;
        RECT 73.430 177.500 73.740 177.550 ;
        RECT 69.470 177.070 69.800 177.170 ;
        RECT 70.640 177.070 70.920 177.240 ;
        RECT 69.470 176.850 70.920 177.070 ;
        RECT 69.470 176.710 69.800 176.850 ;
        RECT 70.640 176.720 70.920 176.850 ;
        RECT 63.270 175.650 63.750 176.320 ;
        RECT 73.960 176.250 74.440 176.410 ;
        RECT 73.960 175.800 74.470 176.250 ;
        RECT 63.290 162.090 63.710 175.650 ;
        RECT 63.290 161.420 63.880 162.090 ;
        RECT 69.980 162.050 70.570 162.260 ;
        RECT 74.030 162.050 74.470 175.800 ;
        RECT 69.980 161.690 74.470 162.050 ;
        RECT 69.980 161.550 70.570 161.690 ;
        RECT 63.290 161.380 63.710 161.420 ;
        RECT 78.580 155.020 79.100 177.550 ;
        RECT 81.780 177.470 87.140 177.690 ;
        RECT 90.120 177.470 90.500 177.560 ;
        RECT 81.780 177.260 90.500 177.470 ;
        RECT 81.780 177.200 87.140 177.260 ;
        RECT 81.780 176.700 82.830 177.200 ;
        RECT 86.690 177.130 87.140 177.200 ;
        RECT 90.120 177.120 90.500 177.260 ;
        RECT 91.340 177.120 91.620 180.470 ;
        RECT 92.490 180.630 92.760 180.790 ;
        RECT 94.140 180.640 94.400 180.780 ;
        RECT 105.700 180.640 106.200 183.760 ;
        RECT 121.190 183.490 121.810 185.000 ;
        RECT 109.320 181.640 109.690 181.810 ;
        RECT 110.550 181.640 110.830 181.750 ;
        RECT 109.320 181.430 110.830 181.640 ;
        RECT 109.320 181.240 109.690 181.430 ;
        RECT 110.550 181.340 110.830 181.430 ;
        RECT 111.560 181.630 111.960 181.800 ;
        RECT 112.860 181.630 113.130 181.770 ;
        RECT 111.560 181.470 113.130 181.630 ;
        RECT 111.560 181.360 111.960 181.470 ;
        RECT 112.860 181.340 113.130 181.470 ;
        RECT 109.920 181.030 110.300 181.170 ;
        RECT 111.130 181.030 111.400 181.180 ;
        RECT 109.920 180.800 111.400 181.030 ;
        RECT 109.920 180.660 110.300 180.800 ;
        RECT 94.140 180.630 106.200 180.640 ;
        RECT 92.490 180.390 106.200 180.630 ;
        RECT 92.490 180.300 92.760 180.390 ;
        RECT 94.140 180.280 106.200 180.390 ;
        RECT 94.140 180.260 105.870 180.280 ;
        RECT 102.990 178.060 104.150 178.080 ;
        RECT 106.470 178.060 106.920 178.100 ;
        RECT 102.990 177.800 106.920 178.060 ;
        RECT 109.900 177.800 110.280 177.890 ;
        RECT 102.990 177.590 110.280 177.800 ;
        RECT 92.380 177.310 92.880 177.530 ;
        RECT 102.990 177.460 106.920 177.590 ;
        RECT 102.990 177.440 106.770 177.460 ;
        RECT 109.900 177.450 110.280 177.590 ;
        RECT 111.120 177.450 111.400 180.800 ;
        RECT 112.270 180.960 112.540 181.120 ;
        RECT 113.920 180.960 114.180 181.110 ;
        RECT 112.270 180.950 114.180 180.960 ;
        RECT 121.180 180.950 121.810 183.490 ;
        RECT 112.270 180.860 121.910 180.950 ;
        RECT 126.000 180.860 126.540 181.090 ;
        RECT 127.190 180.860 127.510 181.020 ;
        RECT 128.940 180.860 129.370 181.070 ;
        RECT 112.270 180.810 126.780 180.860 ;
        RECT 127.190 180.810 129.370 180.860 ;
        RECT 112.270 180.720 129.370 180.810 ;
        RECT 112.270 180.630 112.540 180.720 ;
        RECT 113.920 180.650 129.370 180.720 ;
        RECT 113.920 180.590 114.180 180.650 ;
        RECT 121.140 180.620 129.370 180.650 ;
        RECT 121.140 180.580 126.780 180.620 ;
        RECT 127.190 180.590 129.370 180.620 ;
        RECT 126.000 180.510 126.540 180.580 ;
        RECT 127.190 180.450 127.510 180.590 ;
        RECT 128.940 180.460 129.370 180.590 ;
        RECT 131.300 180.760 131.760 185.100 ;
        RECT 137.310 180.760 138.470 181.060 ;
        RECT 128.360 179.950 128.660 180.210 ;
        RECT 129.570 179.950 129.870 180.230 ;
        RECT 131.300 180.100 138.470 180.760 ;
        RECT 131.300 180.080 131.760 180.100 ;
        RECT 131.300 180.030 131.710 180.080 ;
        RECT 128.360 179.710 129.870 179.950 ;
        RECT 137.310 179.940 138.470 180.100 ;
        RECT 128.360 179.520 128.660 179.710 ;
        RECT 129.570 179.540 129.870 179.710 ;
        RECT 143.400 178.630 143.760 186.460 ;
        RECT 140.650 178.010 141.040 178.160 ;
        RECT 143.400 178.070 143.810 178.630 ;
        RECT 141.810 178.010 143.810 178.070 ;
        RECT 112.160 177.640 112.660 177.860 ;
        RECT 140.650 177.810 143.810 178.010 ;
        RECT 140.650 177.790 143.730 177.810 ;
        RECT 140.650 177.770 142.230 177.790 ;
        RECT 115.630 177.640 115.940 177.710 ;
        RECT 112.160 177.570 115.940 177.640 ;
        RECT 121.170 177.650 122.010 177.660 ;
        RECT 118.850 177.570 119.370 177.610 ;
        RECT 95.850 177.310 96.160 177.380 ;
        RECT 92.380 177.270 96.160 177.310 ;
        RECT 101.170 177.270 101.850 177.340 ;
        RECT 81.830 161.090 82.830 176.700 ;
        RECT 89.440 176.910 89.930 176.950 ;
        RECT 90.700 176.910 91.030 177.000 ;
        RECT 89.440 176.650 91.120 176.910 ;
        RECT 89.440 176.630 91.030 176.650 ;
        RECT 89.440 176.400 89.930 176.630 ;
        RECT 90.700 176.540 91.030 176.630 ;
        RECT 91.340 176.530 91.640 177.120 ;
        RECT 92.380 176.900 101.850 177.270 ;
        RECT 92.380 176.780 92.880 176.900 ;
        RECT 95.850 176.820 96.160 176.900 ;
        RECT 91.890 176.390 92.220 176.490 ;
        RECT 93.060 176.390 93.340 176.560 ;
        RECT 91.890 176.170 93.340 176.390 ;
        RECT 91.890 176.030 92.220 176.170 ;
        RECT 93.060 176.040 93.340 176.170 ;
        RECT 85.590 175.440 86.160 175.630 ;
        RECT 85.590 174.960 86.230 175.440 ;
        RECT 96.390 175.040 97.020 175.760 ;
        RECT 85.730 162.700 86.230 174.960 ;
        RECT 92.620 162.960 93.250 163.020 ;
        RECT 96.470 163.000 96.970 175.040 ;
        RECT 95.370 162.960 96.970 163.000 ;
        RECT 85.730 162.030 86.300 162.700 ;
        RECT 92.620 162.410 96.970 162.960 ;
        RECT 92.620 162.300 93.250 162.410 ;
        RECT 95.370 162.340 96.970 162.410 ;
        RECT 81.670 159.510 82.900 161.090 ;
        RECT 81.830 159.450 82.830 159.510 ;
        RECT 101.170 155.020 101.850 176.900 ;
        RECT 102.990 166.740 104.150 177.440 ;
        RECT 109.220 177.240 109.710 177.280 ;
        RECT 110.480 177.240 110.810 177.330 ;
        RECT 109.220 176.980 110.900 177.240 ;
        RECT 109.220 176.960 110.810 176.980 ;
        RECT 109.220 176.730 109.710 176.960 ;
        RECT 110.480 176.870 110.810 176.960 ;
        RECT 111.120 176.860 111.420 177.450 ;
        RECT 112.160 177.230 119.370 177.570 ;
        RECT 112.160 177.110 112.660 177.230 ;
        RECT 115.560 177.190 119.370 177.230 ;
        RECT 115.630 177.150 115.940 177.190 ;
        RECT 111.670 176.720 112.000 176.820 ;
        RECT 112.840 176.720 113.120 176.890 ;
        RECT 111.670 176.500 113.120 176.720 ;
        RECT 111.670 176.360 112.000 176.500 ;
        RECT 112.840 176.370 113.120 176.500 ;
        RECT 105.300 175.860 105.880 175.930 ;
        RECT 102.900 162.750 104.250 166.740 ;
        RECT 105.300 163.360 105.940 175.860 ;
        RECT 116.130 164.410 116.740 176.080 ;
        RECT 116.130 163.550 116.690 164.410 ;
        RECT 103.040 162.220 104.070 162.750 ;
        RECT 105.180 162.420 107.310 163.360 ;
        RECT 113.570 163.020 116.690 163.550 ;
        RECT 113.570 162.830 114.050 163.020 ;
        RECT 78.490 153.720 102.460 155.020 ;
        RECT 60.140 153.150 73.500 153.190 ;
        RECT 60.140 152.970 73.780 153.150 ;
        RECT 81.480 152.970 82.710 153.130 ;
        RECT 93.240 152.970 93.880 153.050 ;
        RECT 97.420 152.970 98.560 153.400 ;
        RECT 101.700 153.390 102.460 153.720 ;
        RECT 60.140 152.300 98.560 152.970 ;
        RECT 60.140 152.270 70.970 152.300 ;
        RECT 72.920 152.050 98.560 152.300 ;
        RECT 81.480 151.550 82.710 152.050 ;
        RECT 92.990 145.940 94.070 152.050 ;
        RECT 97.420 151.640 98.560 152.050 ;
        RECT 101.550 152.730 102.690 153.390 ;
        RECT 118.850 152.730 119.370 177.190 ;
        RECT 121.170 177.560 125.340 177.650 ;
        RECT 140.650 177.570 141.040 177.770 ;
        RECT 121.170 177.510 127.880 177.560 ;
        RECT 121.170 177.220 127.890 177.510 ;
        RECT 142.080 177.480 142.550 177.520 ;
        RECT 141.790 177.470 142.550 177.480 ;
        RECT 135.890 177.260 136.240 177.270 ;
        RECT 121.170 176.920 125.340 177.220 ;
        RECT 121.170 157.440 122.010 176.920 ;
        RECT 127.670 175.260 127.890 177.220 ;
        RECT 132.020 177.210 136.240 177.260 ;
        RECT 129.970 176.960 136.240 177.210 ;
        RECT 129.970 176.920 132.350 176.960 ;
        RECT 124.480 166.420 125.220 174.560 ;
        RECT 127.530 174.530 128.040 175.260 ;
        RECT 129.980 175.150 130.180 176.920 ;
        RECT 132.020 176.860 132.350 176.920 ;
        RECT 129.910 174.580 130.300 175.150 ;
        RECT 127.000 173.850 127.360 174.000 ;
        RECT 128.190 173.850 128.550 174.020 ;
        RECT 127.000 173.610 128.550 173.850 ;
        RECT 127.000 173.460 127.360 173.610 ;
        RECT 128.190 173.480 128.550 173.610 ;
        RECT 129.330 173.880 129.690 174.090 ;
        RECT 130.500 173.880 130.860 174.090 ;
        RECT 129.330 173.620 130.860 173.880 ;
        RECT 132.780 173.760 133.420 174.440 ;
        RECT 129.330 173.440 129.690 173.620 ;
        RECT 130.500 173.440 130.860 173.620 ;
        RECT 123.940 166.020 125.220 166.420 ;
        RECT 123.940 163.130 124.680 166.020 ;
        RECT 123.940 162.450 124.770 163.130 ;
        RECT 130.930 163.110 131.570 163.280 ;
        RECT 132.930 163.110 133.370 173.760 ;
        RECT 135.890 171.440 136.240 176.960 ;
        RECT 139.820 177.100 140.480 177.470 ;
        RECT 141.200 177.100 142.550 177.470 ;
        RECT 139.820 176.740 142.550 177.100 ;
        RECT 139.820 176.560 140.480 176.740 ;
        RECT 141.200 176.560 142.550 176.740 ;
        RECT 135.880 170.980 136.240 171.440 ;
        RECT 135.880 166.480 136.230 170.980 ;
        RECT 130.930 162.780 133.370 163.110 ;
        RECT 130.930 162.600 131.570 162.780 ;
        RECT 124.100 162.180 124.770 162.450 ;
        RECT 121.170 155.810 122.310 157.440 ;
        RECT 135.500 154.070 136.590 166.480 ;
        RECT 142.080 165.370 142.550 176.560 ;
        RECT 140.350 165.110 140.900 165.250 ;
        RECT 141.660 165.110 142.550 165.370 ;
        RECT 140.350 164.900 142.550 165.110 ;
        RECT 140.350 164.680 142.210 164.900 ;
        RECT 140.350 164.500 140.900 164.680 ;
        RECT 141.660 164.620 142.210 164.680 ;
        RECT 141.110 163.630 141.400 163.800 ;
        RECT 143.200 163.630 143.480 163.640 ;
        RECT 141.110 163.390 143.480 163.630 ;
        RECT 141.110 163.270 141.400 163.390 ;
        RECT 130.400 152.730 131.700 153.100 ;
        RECT 135.500 152.730 136.550 154.070 ;
        RECT 143.200 153.160 143.480 163.390 ;
        RECT 101.550 152.020 136.550 152.730 ;
        RECT 101.550 151.630 102.690 152.020 ;
        RECT 121.320 149.890 122.560 150.980 ;
        RECT 130.400 150.910 131.700 152.020 ;
        RECT 135.500 151.970 136.550 152.020 ;
        RECT 143.150 152.330 143.550 153.160 ;
        RECT 121.560 145.940 122.250 149.890 ;
        RECT 92.990 145.880 122.400 145.940 ;
        RECT 143.150 145.880 143.520 152.330 ;
        RECT 92.990 145.470 143.520 145.880 ;
        RECT 92.970 144.840 143.520 145.470 ;
        RECT 92.970 144.710 122.400 144.840 ;
        RECT 92.970 142.600 94.890 144.710 ;
        RECT 92.970 142.000 94.980 142.600 ;
        RECT 92.940 140.470 94.980 142.000 ;
        RECT 93.190 139.900 94.980 140.470 ;
        RECT 130.170 139.480 131.960 141.490 ;
        RECT 100.810 113.120 101.310 113.200 ;
        RECT 68.090 112.880 68.590 112.960 ;
        RECT 100.810 112.930 107.800 113.120 ;
        RECT 100.810 112.920 107.310 112.930 ;
        RECT 68.090 112.690 75.080 112.880 ;
        RECT 100.810 112.800 101.310 112.920 ;
        RECT 68.090 112.680 74.590 112.690 ;
        RECT 68.090 112.560 68.590 112.680 ;
        RECT 74.760 112.050 75.080 112.690 ;
        RECT 107.480 112.290 107.800 112.930 ;
        RECT 74.680 111.420 75.290 112.050 ;
        RECT 107.400 111.660 108.010 112.290 ;
        RECT 56.680 101.950 58.750 104.950 ;
        RECT 94.130 104.790 95.030 105.350 ;
        RECT 105.920 104.790 106.480 105.020 ;
        RECT 73.030 104.530 73.660 104.740 ;
        RECT 79.400 104.530 79.910 104.560 ;
        RECT 73.030 104.110 79.910 104.530 ;
        RECT 94.130 104.430 106.480 104.790 ;
        RECT 94.130 104.200 95.030 104.430 ;
        RECT 105.920 104.200 106.480 104.430 ;
        RECT 73.030 104.060 73.660 104.110 ;
        RECT 79.400 103.680 79.910 104.110 ;
        RECT 57.510 74.150 58.160 101.950 ;
        RECT 79.400 100.370 79.920 103.680 ;
        RECT 71.950 99.250 72.360 99.420 ;
        RECT 73.180 99.250 73.480 99.330 ;
        RECT 71.950 99.020 73.480 99.250 ;
        RECT 71.950 98.970 72.360 99.020 ;
        RECT 73.180 98.890 73.480 99.020 ;
        RECT 62.550 97.790 63.520 98.770 ;
        RECT 79.380 94.340 79.920 100.370 ;
        RECT 104.670 99.490 105.080 99.660 ;
        RECT 105.900 99.490 106.200 99.570 ;
        RECT 104.670 99.260 106.200 99.490 ;
        RECT 104.670 99.210 105.080 99.260 ;
        RECT 105.900 99.130 106.200 99.260 ;
        RECT 95.310 98.010 96.090 98.770 ;
        RECT 79.380 93.100 79.900 94.340 ;
        RECT 79.100 91.660 80.230 93.100 ;
        RECT 99.460 87.020 99.960 87.100 ;
        RECT 99.460 86.830 106.450 87.020 ;
        RECT 99.460 86.820 105.960 86.830 ;
        RECT 99.460 86.700 99.960 86.820 ;
        RECT 106.130 86.190 106.450 86.830 ;
        RECT 106.050 85.560 106.660 86.190 ;
        RECT 67.810 84.500 68.310 84.580 ;
        RECT 67.810 84.310 74.800 84.500 ;
        RECT 67.810 84.300 74.310 84.310 ;
        RECT 67.810 84.180 68.310 84.300 ;
        RECT 74.480 83.670 74.800 84.310 ;
        RECT 74.400 83.040 75.010 83.670 ;
        RECT 104.450 78.780 105.030 78.910 ;
        RECT 91.230 78.180 105.030 78.780 ;
        RECT 91.230 78.020 93.540 78.180 ;
        RECT 91.390 77.720 92.190 78.020 ;
        RECT 85.570 76.460 86.690 76.540 ;
        RECT 72.730 75.760 86.740 76.460 ;
        RECT 72.730 75.710 73.380 75.760 ;
        RECT 61.240 74.150 62.010 74.560 ;
        RECT 57.510 73.740 62.180 74.150 ;
        RECT 61.240 73.570 62.010 73.740 ;
        RECT 71.670 70.870 72.080 71.040 ;
        RECT 72.900 70.870 73.200 70.950 ;
        RECT 71.670 70.640 73.200 70.870 ;
        RECT 71.670 70.590 72.080 70.640 ;
        RECT 72.900 70.510 73.200 70.640 ;
        RECT 85.570 63.390 86.690 75.760 ;
        RECT 91.300 72.060 92.190 77.720 ;
        RECT 99.280 76.770 100.070 76.900 ;
        RECT 92.940 76.010 100.070 76.770 ;
        RECT 92.940 75.930 99.950 76.010 ;
        RECT 91.300 67.350 92.090 72.060 ;
        RECT 92.980 69.180 93.690 75.930 ;
        RECT 103.320 73.390 103.730 73.560 ;
        RECT 104.550 73.390 104.850 73.470 ;
        RECT 103.320 73.160 104.850 73.390 ;
        RECT 103.320 73.110 103.730 73.160 ;
        RECT 104.550 73.030 104.850 73.160 ;
        RECT 92.980 69.130 93.520 69.180 ;
        RECT 91.300 66.620 92.190 67.350 ;
        RECT 91.390 63.600 92.190 66.620 ;
        RECT 85.430 61.890 86.920 63.390 ;
        RECT 91.030 62.350 92.420 63.600 ;
        RECT 73.070 58.570 73.490 58.800 ;
        RECT 76.150 58.570 76.570 58.800 ;
        RECT 73.070 58.340 76.580 58.570 ;
        RECT 73.070 58.280 73.490 58.340 ;
        RECT 76.150 58.280 76.570 58.340 ;
        RECT 87.480 57.410 87.900 57.640 ;
        RECT 90.560 57.410 90.980 57.640 ;
        RECT 87.480 57.180 90.990 57.410 ;
        RECT 87.480 57.120 87.900 57.180 ;
        RECT 90.560 57.120 90.980 57.180 ;
        RECT 73.150 56.600 73.500 56.650 ;
        RECT 73.090 56.590 73.980 56.600 ;
        RECT 76.160 56.590 76.560 56.720 ;
        RECT 73.090 56.580 74.250 56.590 ;
        RECT 75.690 56.580 76.560 56.590 ;
        RECT 73.090 56.340 76.560 56.580 ;
        RECT 73.090 56.330 73.980 56.340 ;
        RECT 73.150 56.250 73.500 56.330 ;
        RECT 75.690 56.300 76.560 56.340 ;
        RECT 76.160 56.240 76.560 56.300 ;
        RECT 87.560 55.440 87.910 55.490 ;
        RECT 87.500 55.430 88.390 55.440 ;
        RECT 90.570 55.430 90.970 55.560 ;
        RECT 87.500 55.420 88.660 55.430 ;
        RECT 90.100 55.420 90.970 55.430 ;
        RECT 87.500 55.180 90.970 55.420 ;
        RECT 87.500 55.170 88.390 55.180 ;
        RECT 87.560 55.090 87.910 55.170 ;
        RECT 90.100 55.140 90.970 55.180 ;
        RECT 90.570 55.080 90.970 55.140 ;
        RECT 38.920 47.980 41.000 49.290 ;
        RECT 38.920 47.910 56.830 47.980 ;
        RECT 38.920 47.640 83.750 47.910 ;
        RECT 38.920 47.230 83.810 47.640 ;
        RECT 39.050 47.090 83.810 47.230 ;
        RECT 39.550 47.030 56.830 47.090 ;
        RECT 82.610 46.410 83.810 47.090 ;
      LAYER met3 ;
        RECT 94.480 210.590 95.160 210.645 ;
        RECT 98.260 210.590 98.780 210.635 ;
        RECT 94.480 210.540 98.780 210.590 ;
        RECT 99.290 210.540 100.000 210.665 ;
        RECT 103.110 210.540 103.820 210.715 ;
        RECT 94.480 210.290 103.820 210.540 ;
        RECT 94.480 210.045 95.160 210.290 ;
        RECT 98.200 210.220 103.820 210.290 ;
        RECT 98.260 210.095 98.780 210.220 ;
        RECT 99.290 209.985 100.000 210.220 ;
        RECT 103.110 210.035 103.820 210.220 ;
        RECT 94.470 206.760 95.060 206.925 ;
        RECT 98.270 206.760 98.860 206.935 ;
        RECT 99.410 206.760 100.000 206.995 ;
        RECT 103.170 206.760 103.760 206.955 ;
        RECT 94.470 206.460 103.760 206.760 ;
        RECT 94.470 206.385 95.060 206.460 ;
        RECT 98.270 206.395 98.860 206.460 ;
        RECT 99.410 206.455 100.000 206.460 ;
        RECT 103.170 206.415 103.760 206.460 ;
        RECT 94.440 203.170 95.050 203.315 ;
        RECT 98.270 203.170 98.880 203.315 ;
        RECT 99.380 203.170 99.970 203.345 ;
        RECT 103.180 203.170 103.770 203.375 ;
        RECT 94.440 202.860 103.770 203.170 ;
        RECT 94.440 202.705 95.050 202.860 ;
        RECT 98.270 202.705 98.880 202.860 ;
        RECT 99.380 202.695 99.970 202.860 ;
        RECT 103.180 202.725 103.770 202.860 ;
        RECT 62.500 98.650 63.570 98.745 ;
        RECT 95.260 98.650 96.140 98.745 ;
        RECT 62.500 98.035 96.140 98.650 ;
        RECT 62.500 97.840 96.120 98.035 ;
        RECT 62.500 97.815 63.570 97.840 ;
  END
END tt_um_subdiduntil2_mixed_signal_classifier
END LIBRARY

