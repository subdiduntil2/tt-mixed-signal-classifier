magic
tech sky130A
magscale 1 2
timestamp 1755904430
<< viali >>
rect 30142 5742 30184 5818
rect 12014 4812 12066 4814
rect 11996 4666 12066 4812
rect 30230 3142 30266 3196
rect 11944 974 11978 1014
rect 22040 -412 22084 -344
rect 22854 -416 22898 -348
<< metal1 >>
rect 11818 7674 12018 7786
rect 11818 7586 12030 7674
rect 11924 7170 12030 7586
rect 11926 6968 12030 7170
rect 13576 7338 13736 7346
rect 15194 7338 16116 7344
rect 13576 7330 16116 7338
rect 17040 7330 17116 7332
rect 13576 7260 17116 7330
rect 13576 7214 16116 7260
rect 13332 6968 13342 6986
rect 11926 6836 13342 6968
rect 11926 6768 12030 6836
rect 13332 6828 13342 6836
rect 13458 6828 13468 6986
rect 11924 6458 12030 6768
rect 13576 6660 13736 7214
rect 17040 7202 17116 7260
rect 20478 7202 24584 7204
rect 17040 7182 28606 7202
rect 17040 7176 28630 7182
rect 17040 7096 28450 7176
rect 20478 7078 28450 7096
rect 24146 7042 28450 7078
rect 24146 7040 24590 7042
rect 15946 6912 15968 6964
rect 15958 6850 15968 6912
rect 16126 6936 16144 6964
rect 16126 6850 16136 6936
rect 24146 6908 24178 7040
rect 28440 7032 28450 7042
rect 28608 7042 28630 7176
rect 28608 7032 28618 7042
rect 20470 6728 20480 6808
rect 20588 6728 20598 6808
rect 24408 6770 24418 6866
rect 24536 6770 24546 6866
rect 11456 6250 11466 6330
rect 11548 6250 11558 6330
rect 11464 6154 11542 6250
rect 11464 6152 11632 6154
rect 11464 6126 11876 6152
rect 11464 6080 11542 6126
rect 11586 6122 11876 6126
rect 11926 6082 12030 6458
rect 13562 6368 13738 6660
rect 13562 6224 13594 6368
rect 13710 6224 13738 6368
rect 13562 6212 13738 6224
rect 27422 6114 27432 6210
rect 27540 6114 27550 6210
rect 28528 6128 28620 6168
rect 11464 5944 11550 6080
rect 11920 6076 12030 6082
rect 11632 6002 11642 6068
rect 11696 6002 11706 6068
rect 11744 5992 11754 6072
rect 11830 5992 11840 6072
rect 11890 5986 11900 6076
rect 11962 5986 12030 6076
rect 17422 5992 17438 6100
rect 11920 5966 12030 5986
rect 11456 5934 11600 5944
rect 11714 5934 11750 5940
rect 11456 5916 11886 5934
rect 11464 5840 11550 5916
rect 11596 5904 11886 5916
rect 11714 5840 11750 5904
rect 11464 5812 11882 5840
rect 11464 5624 11550 5812
rect 11592 5810 11882 5812
rect 11714 5806 11750 5810
rect 11920 5758 12006 5966
rect 25746 5938 27174 6054
rect 28482 6018 28492 6128
rect 28574 6094 28620 6128
rect 28574 6062 28610 6094
rect 28574 6056 28624 6062
rect 28574 6018 28584 6056
rect 29684 6000 29694 6204
rect 29926 6168 29936 6204
rect 30120 6168 31032 6172
rect 29926 6056 31196 6168
rect 29926 6000 29936 6056
rect 11630 5686 11640 5752
rect 11694 5686 11704 5752
rect 11744 5674 11754 5754
rect 11830 5674 11840 5754
rect 11892 5668 11902 5758
rect 11964 5668 12006 5758
rect 11464 5622 11616 5624
rect 11464 5592 11884 5622
rect 11464 5514 11550 5592
rect 11714 5516 11750 5592
rect 11920 5540 12006 5668
rect 11920 5526 12020 5540
rect 11920 5522 12034 5526
rect 11756 5516 11878 5518
rect 11464 5482 11598 5514
rect 11624 5486 11878 5516
rect 11756 5482 11878 5486
rect 11922 5486 12034 5522
rect 11922 5482 12020 5486
rect 11464 5300 11550 5482
rect 11920 5478 12020 5482
rect 11640 5362 11650 5428
rect 11704 5362 11714 5428
rect 11752 5348 11762 5444
rect 11838 5348 11848 5444
rect 11920 5438 12006 5478
rect 11884 5348 11894 5438
rect 11956 5348 12006 5438
rect 11464 5298 11596 5300
rect 11712 5298 11748 5302
rect 11464 5268 11872 5298
rect 11464 5190 11550 5268
rect 11712 5192 11748 5268
rect 11596 5190 11886 5192
rect 11464 5162 11886 5190
rect 11464 5158 11604 5162
rect 11464 4982 11550 5158
rect 11636 5040 11646 5106
rect 11700 5040 11710 5106
rect 11748 5030 11758 5126
rect 11834 5030 11844 5126
rect 11920 5116 12006 5348
rect 14876 5142 14886 5256
rect 14982 5142 14992 5256
rect 17014 5172 17024 5274
rect 17120 5172 17130 5274
rect 11878 5026 11888 5116
rect 11950 5026 12006 5116
rect 11464 4980 11600 4982
rect 11464 4950 11882 4980
rect 11464 4874 11550 4950
rect 11720 4876 11756 4950
rect 11614 4874 11886 4876
rect 11464 4846 11886 4874
rect 11920 4846 12006 5026
rect 19340 5004 19350 5118
rect 19464 5004 19474 5118
rect 21500 5020 21510 5144
rect 21636 5020 21646 5144
rect 23282 5058 23292 5178
rect 23408 5058 23418 5178
rect 25462 5068 25472 5192
rect 25568 5068 25578 5192
rect 11464 4842 11622 4846
rect 11720 4844 11756 4846
rect 11464 4664 11550 4842
rect 11920 4814 17442 4846
rect 11920 4812 12014 4814
rect 11640 4720 11650 4786
rect 11704 4720 11714 4786
rect 11756 4706 11766 4802
rect 11842 4706 11852 4802
rect 11920 4800 11996 4812
rect 11882 4710 11892 4800
rect 11954 4710 11996 4800
rect 11920 4666 11996 4710
rect 12066 4718 17442 4814
rect 25850 4748 25938 5938
rect 28414 5818 30200 5842
rect 28414 5742 30142 5818
rect 30184 5742 30200 5818
rect 28414 5714 30200 5742
rect 30372 5716 30442 6056
rect 28414 5708 28786 5714
rect 27134 4806 27144 4902
rect 27276 4806 27286 4902
rect 28778 4764 28788 4880
rect 28916 4764 28926 4880
rect 12066 4710 19944 4718
rect 12066 4704 21768 4710
rect 12066 4666 24436 4704
rect 11464 4632 11608 4664
rect 11718 4658 11754 4662
rect 11464 4556 11550 4632
rect 11610 4628 11884 4658
rect 11718 4560 11754 4628
rect 11920 4626 24436 4666
rect 11604 4556 11884 4560
rect 11464 4530 11884 4556
rect 11464 4524 11626 4530
rect 11718 4528 11754 4530
rect 11464 4348 11550 4524
rect 11636 4398 11646 4464
rect 11700 4398 11710 4464
rect 11744 4386 11754 4482
rect 11830 4386 11840 4482
rect 11920 4476 12006 4626
rect 11878 4386 11888 4476
rect 11950 4386 12006 4476
rect 11464 4346 11624 4348
rect 11464 4316 11876 4346
rect 11464 4242 11550 4316
rect 11464 4236 11614 4242
rect 11714 4236 11750 4316
rect 11464 4210 11848 4236
rect 11464 4166 11554 4210
rect 11608 4198 11848 4210
rect 11462 4068 11554 4166
rect 11628 4080 11638 4140
rect 11694 4080 11704 4140
rect 11748 4074 11758 4160
rect 11838 4074 11848 4160
rect 11920 4148 12006 4386
rect 11880 4078 11890 4148
rect 11944 4078 12006 4148
rect 11464 4022 11554 4068
rect 11464 3992 11878 4022
rect 11464 3986 11588 3992
rect 11464 3916 11550 3986
rect 11464 3914 11604 3916
rect 11712 3914 11748 3992
rect 11464 3884 11882 3914
rect 11464 3702 11550 3884
rect 11920 3840 12006 4078
rect 11632 3762 11642 3828
rect 11696 3762 11706 3828
rect 11752 3750 11762 3830
rect 11838 3750 11848 3830
rect 11886 3750 11896 3840
rect 11958 3750 12006 3840
rect 11464 3670 11604 3702
rect 11608 3678 11884 3708
rect 11464 3594 11550 3670
rect 11716 3602 11752 3678
rect 11596 3594 11886 3602
rect 11464 3572 11886 3594
rect 11464 3562 11604 3572
rect 11716 3564 11752 3572
rect 11464 3382 11550 3562
rect 11920 3522 12006 3750
rect 11632 3446 11642 3512
rect 11696 3446 11706 3512
rect 11744 3434 11754 3514
rect 11830 3434 11840 3514
rect 11878 3432 11888 3522
rect 11950 3432 12006 3522
rect 11464 3374 11606 3382
rect 11464 3350 11882 3374
rect 11464 3278 11550 3350
rect 11592 3344 11882 3350
rect 11464 3270 11608 3278
rect 11712 3270 11744 3344
rect 11464 3246 11882 3270
rect 11464 3166 11550 3246
rect 11592 3240 11882 3246
rect 11920 3200 12006 3432
rect 11462 3064 11556 3166
rect 11628 3120 11638 3186
rect 11692 3120 11702 3186
rect 11750 3118 11760 3198
rect 11836 3118 11846 3198
rect 11884 3110 11894 3200
rect 11956 3124 12006 3200
rect 11956 3110 11966 3124
rect 11462 3062 11602 3064
rect 11462 3032 11878 3062
rect 11462 3030 11556 3032
rect 12432 2246 12752 4626
rect 15138 2746 15342 4626
rect 17172 4570 24436 4626
rect 25660 4604 26112 4748
rect 17172 4566 23510 4570
rect 17172 4564 19944 4566
rect 19636 2922 19846 4564
rect 21664 4550 23510 4566
rect 23804 4550 24436 4570
rect 23860 2998 23998 4550
rect 25994 3036 26112 4604
rect 29798 3208 29920 5714
rect 30326 5684 30472 5716
rect 30352 5526 30362 5624
rect 30440 5526 30450 5624
rect 31084 5562 31192 6056
rect 31078 5530 31192 5562
rect 30186 5324 30196 5486
rect 30328 5324 30338 5486
rect 30462 5324 30472 5486
rect 30604 5324 30614 5486
rect 30320 5050 30466 5082
rect 30398 4762 30446 5050
rect 31078 4766 31190 5530
rect 30870 4762 31190 4766
rect 30398 4696 31190 4762
rect 30398 4694 31176 4696
rect 30398 4692 30890 4694
rect 30398 3504 30446 4692
rect 30394 3458 31028 3504
rect 29798 3196 30292 3208
rect 29798 3142 30230 3196
rect 30266 3142 30292 3196
rect 30398 3160 30446 3458
rect 30398 3150 30572 3160
rect 29798 3122 30292 3142
rect 30426 3128 30572 3150
rect 25994 2954 27454 3036
rect 19772 2890 19846 2922
rect 30292 2912 30302 3042
rect 30412 2912 30422 3042
rect 30554 2936 30564 3066
rect 30674 2936 30684 3066
rect 19024 2508 19224 2598
rect 19368 2508 19378 2532
rect 14492 2382 14692 2446
rect 14902 2382 14912 2410
rect 14492 2296 14912 2382
rect 15008 2296 15018 2410
rect 16218 2322 16228 2444
rect 16346 2322 16356 2444
rect 19024 2420 19378 2508
rect 14492 2280 14958 2296
rect 14492 2246 14692 2280
rect 11856 2242 12756 2246
rect 11852 2216 12756 2242
rect 11852 2100 11880 2216
rect 11614 2062 11884 2100
rect 11514 1976 11524 1990
rect 11452 1894 11524 1976
rect 11610 1894 11620 1990
rect 11748 1902 11758 1998
rect 11844 1902 11854 1998
rect 11452 1652 11552 1894
rect 11630 1734 11640 1830
rect 11726 1734 11736 1830
rect 11868 1734 11878 1830
rect 11964 1734 11974 1830
rect 11436 1556 11552 1652
rect 11622 1630 11892 1652
rect 12432 1630 12752 2216
rect 18540 2210 18812 2420
rect 19024 2398 19224 2420
rect 19368 2418 19378 2420
rect 19492 2508 19502 2532
rect 19492 2420 19522 2508
rect 20746 2472 20756 2596
rect 20882 2472 20892 2596
rect 22830 2456 22840 2700
rect 23046 2456 23056 2700
rect 23528 2642 23712 2678
rect 23528 2618 23556 2642
rect 23310 2528 23556 2618
rect 19492 2418 19502 2420
rect 11452 1440 11552 1556
rect 11600 1516 12752 1630
rect 11620 1510 11890 1516
rect 11452 1360 11528 1440
rect 11610 1360 11620 1440
rect 11762 1372 11772 1452
rect 11854 1372 11864 1452
rect 11452 1350 11552 1360
rect 11644 1198 11654 1278
rect 11736 1198 11746 1278
rect 11940 1268 12004 1278
rect 11880 1188 11890 1268
rect 11972 1188 12004 1268
rect 11608 1066 11878 1104
rect 11714 922 11776 1066
rect 11932 1014 12004 1188
rect 11932 974 11944 1014
rect 11978 974 12004 1014
rect 11660 790 11670 922
rect 11794 790 11804 922
rect 11932 776 12004 974
rect 12616 934 12750 1516
rect 14958 1080 15112 1932
rect 18540 1914 18566 2210
rect 18812 1914 18822 2210
rect 12596 780 12606 934
rect 12734 914 12750 934
rect 12734 780 12744 914
rect 11902 734 12102 776
rect 14942 734 15114 1080
rect 11902 612 15114 734
rect 18540 618 18812 1914
rect 19800 1292 19908 2092
rect 22890 1782 23016 2456
rect 23324 2194 23416 2528
rect 23546 2522 23556 2528
rect 23672 2596 23712 2642
rect 23672 2522 23682 2596
rect 24936 2578 24946 2702
rect 25042 2578 25052 2702
rect 30444 2666 30454 2752
rect 30512 2666 30522 2752
rect 30936 2690 31024 3458
rect 27042 2582 27052 2618
rect 26874 2570 27052 2582
rect 26838 2500 27052 2570
rect 26838 2222 26906 2500
rect 27042 2448 27052 2500
rect 27186 2448 27196 2618
rect 28408 2532 28418 2648
rect 28546 2532 28556 2648
rect 30936 2534 31016 2690
rect 30524 2532 31016 2534
rect 30422 2500 31016 2532
rect 30524 2488 31016 2500
rect 23280 1994 23480 2194
rect 21772 1750 23016 1782
rect 21762 1672 23016 1750
rect 21762 1622 23010 1672
rect 19800 1158 19934 1292
rect 11902 576 12102 612
rect 14942 -280 15114 612
rect 18518 322 18528 618
rect 18774 420 18812 618
rect 18774 322 18784 420
rect 19808 -216 19934 1158
rect 21762 672 21890 1622
rect 23646 962 23818 2206
rect 26782 2022 26982 2222
rect 26456 1174 26466 1480
rect 26694 1174 26704 1480
rect 23640 764 23818 962
rect 20854 602 21054 638
rect 20854 458 20880 602
rect 21008 572 21054 602
rect 21706 572 21716 672
rect 21008 528 21716 572
rect 21008 458 21054 528
rect 20854 438 21054 458
rect 21706 340 21716 528
rect 21944 340 21954 672
rect 22532 338 22542 670
rect 22770 566 22780 670
rect 23088 566 23288 614
rect 22770 436 23288 566
rect 23640 542 23816 764
rect 23640 468 23818 542
rect 22770 338 22780 436
rect 23088 414 23288 436
rect 18494 -220 22892 -216
rect 23646 -220 23818 468
rect 26536 188 26634 1174
rect 26486 -10 26496 188
rect 26744 -10 26754 188
rect 27146 -120 27318 2118
rect 27146 -186 27310 -120
rect 27070 -208 27310 -186
rect 26980 -220 27310 -208
rect 18494 -280 27310 -220
rect 14942 -344 27310 -280
rect 14942 -412 22040 -344
rect 22084 -348 27310 -344
rect 22084 -412 22854 -348
rect 14942 -416 22854 -412
rect 22898 -416 27310 -348
rect 14942 -508 27310 -416
rect 14942 -526 22892 -508
rect 26980 -514 27310 -508
rect 14942 -532 19370 -526
rect 27070 -528 27310 -514
rect 14942 -538 15114 -532
<< via1 >>
rect 13342 6828 13458 6986
rect 15968 6850 16126 6964
rect 28450 7032 28608 7176
rect 20480 6728 20588 6808
rect 24418 6770 24536 6866
rect 11466 6250 11548 6330
rect 13594 6224 13710 6368
rect 27432 6114 27540 6210
rect 11642 6002 11696 6068
rect 11754 5992 11830 6072
rect 11900 5986 11962 6076
rect 28492 6018 28574 6128
rect 29694 6000 29926 6204
rect 11640 5686 11694 5752
rect 11754 5674 11830 5754
rect 11902 5668 11964 5758
rect 11650 5362 11704 5428
rect 11762 5348 11838 5444
rect 11894 5348 11956 5438
rect 11646 5040 11700 5106
rect 11758 5030 11834 5126
rect 14886 5142 14982 5256
rect 17024 5172 17120 5274
rect 11888 5026 11950 5116
rect 19350 5004 19464 5118
rect 21510 5020 21636 5144
rect 23292 5058 23408 5178
rect 25472 5068 25568 5192
rect 11650 4720 11704 4786
rect 11766 4706 11842 4802
rect 11892 4710 11954 4800
rect 27144 4806 27276 4902
rect 28788 4764 28916 4880
rect 11646 4398 11700 4464
rect 11754 4386 11830 4482
rect 11888 4386 11950 4476
rect 11638 4080 11694 4140
rect 11758 4074 11838 4160
rect 11890 4078 11944 4148
rect 11642 3762 11696 3828
rect 11762 3750 11838 3830
rect 11896 3750 11958 3840
rect 11642 3446 11696 3512
rect 11754 3434 11830 3514
rect 11888 3432 11950 3522
rect 11638 3120 11692 3186
rect 11760 3118 11836 3198
rect 11894 3110 11956 3200
rect 30362 5526 30440 5624
rect 30196 5324 30328 5486
rect 30472 5324 30604 5486
rect 30302 2912 30412 3042
rect 30564 2936 30674 3066
rect 14912 2296 15008 2410
rect 16228 2322 16346 2444
rect 11524 1894 11610 1990
rect 11758 1902 11844 1998
rect 11640 1734 11726 1830
rect 11878 1734 11964 1830
rect 19378 2418 19492 2532
rect 20756 2472 20882 2596
rect 22840 2456 23046 2700
rect 11528 1360 11610 1440
rect 11772 1372 11854 1452
rect 11654 1198 11736 1278
rect 11890 1188 11972 1268
rect 11670 790 11794 922
rect 18566 1914 18812 2210
rect 12606 780 12734 934
rect 23556 2522 23672 2642
rect 24946 2578 25042 2702
rect 30454 2666 30512 2752
rect 27052 2448 27186 2618
rect 28418 2532 28546 2648
rect 18528 322 18774 618
rect 26466 1174 26694 1480
rect 20880 458 21008 602
rect 21716 340 21944 672
rect 22542 338 22770 670
rect 26496 -10 26744 188
<< metal2 >>
rect 30912 7418 30984 7424
rect 26470 7294 30984 7418
rect 26470 7246 26610 7294
rect 26454 7028 26610 7246
rect 28492 7186 28584 7198
rect 26470 7002 26610 7028
rect 28450 7182 28606 7186
rect 28450 7176 28608 7182
rect 28608 7042 28630 7140
rect 28450 7022 28608 7032
rect 13342 6986 13458 6996
rect 15968 6964 16126 6974
rect 13458 6850 15968 6948
rect 16126 6850 16130 6948
rect 24418 6866 24536 6876
rect 13458 6828 16130 6850
rect 13342 6818 13458 6828
rect 20480 6808 20588 6818
rect 19432 6728 20480 6798
rect 20588 6728 20594 6798
rect 19432 6682 20594 6728
rect 23372 6770 24418 6854
rect 24536 6770 24560 6854
rect 23372 6754 24560 6770
rect 13594 6368 13710 6378
rect 11466 6330 11548 6340
rect 11446 6294 11466 6324
rect 13374 6324 13594 6326
rect 11548 6270 13594 6324
rect 11548 6268 11824 6270
rect 11466 6240 11548 6250
rect 11632 6090 11722 6100
rect 11764 6082 11824 6268
rect 13374 6260 13594 6270
rect 13594 6214 13710 6224
rect 16582 6282 17470 6296
rect 19432 6282 19542 6682
rect 16582 6210 19542 6282
rect 17618 6202 19542 6210
rect 19432 6196 19542 6202
rect 23372 6130 23472 6754
rect 26470 6700 26594 7002
rect 26468 6192 26594 6700
rect 27432 6210 27540 6220
rect 25026 6174 26614 6192
rect 25026 6132 27432 6174
rect 11880 6092 11970 6102
rect 11754 6072 11830 6082
rect 11754 5982 11830 5992
rect 21074 6058 23472 6130
rect 26460 6118 27432 6132
rect 27540 6164 27588 6174
rect 27540 6126 27708 6164
rect 28492 6154 28584 7022
rect 29694 6204 29926 6214
rect 28492 6128 29694 6154
rect 27540 6118 27588 6126
rect 27432 6104 27540 6114
rect 21074 6054 23406 6058
rect 28574 6022 29694 6128
rect 28574 6018 28584 6022
rect 28492 6008 28574 6018
rect 29694 5990 29926 6000
rect 11632 5962 11722 5972
rect 11620 5774 11710 5784
rect 11764 5764 11824 5982
rect 11880 5964 11970 5974
rect 11882 5778 11972 5788
rect 11754 5754 11830 5764
rect 11754 5664 11830 5674
rect 11620 5646 11710 5656
rect 11626 5458 11716 5468
rect 11764 5454 11824 5664
rect 11882 5650 11972 5660
rect 30912 5728 30984 7294
rect 14268 5598 15380 5654
rect 30362 5624 30440 5634
rect 22830 5614 23062 5618
rect 14268 5556 14398 5598
rect 11880 5458 11970 5468
rect 11626 5330 11716 5340
rect 11762 5444 11838 5454
rect 11762 5338 11838 5348
rect 11638 5132 11728 5142
rect 11764 5136 11824 5338
rect 11880 5330 11970 5340
rect 11758 5126 11834 5136
rect 11758 5020 11834 5030
rect 11876 5132 11966 5142
rect 11638 5004 11728 5014
rect 11764 4962 11824 5020
rect 11876 5004 11966 5014
rect 11626 4816 11716 4826
rect 11626 4688 11716 4698
rect 11764 4812 11834 4962
rect 11880 4812 11970 4822
rect 11764 4802 11842 4812
rect 11764 4706 11766 4802
rect 11764 4696 11842 4706
rect 11628 4488 11714 4498
rect 11764 4492 11834 4696
rect 11880 4684 11970 4694
rect 11754 4482 11834 4492
rect 11830 4386 11834 4482
rect 11754 4376 11834 4386
rect 11628 4364 11714 4374
rect 11628 4164 11726 4174
rect 11764 4170 11834 4376
rect 11876 4490 11962 4500
rect 11876 4366 11962 4376
rect 11628 4056 11726 4066
rect 11758 4160 11838 4170
rect 11758 4064 11838 4074
rect 11870 4166 11966 4176
rect 11630 3856 11720 3866
rect 11768 3840 11824 4064
rect 11870 4058 11966 4068
rect 11874 3860 11964 3870
rect 11762 3830 11838 3840
rect 11762 3740 11838 3750
rect 11630 3728 11720 3738
rect 11626 3534 11716 3544
rect 11768 3524 11824 3740
rect 11874 3732 11964 3742
rect 11872 3532 11962 3542
rect 11754 3514 11830 3524
rect 11754 3424 11830 3434
rect 11626 3406 11716 3416
rect 11618 3214 11708 3224
rect 11768 3208 11824 3424
rect 11872 3404 11962 3414
rect 11880 3212 11970 3222
rect 11760 3198 11836 3208
rect 11760 3108 11836 3118
rect 11618 3086 11708 3096
rect 11776 2008 11824 3108
rect 11880 3084 11970 3094
rect 11524 1990 11610 2000
rect 11758 1998 11844 2008
rect 11610 1920 11758 1978
rect 11524 1884 11610 1894
rect 11758 1892 11844 1902
rect 11640 1830 11726 1840
rect 11878 1830 11964 1840
rect 11726 1762 11878 1820
rect 11640 1724 11726 1734
rect 11964 1734 12014 1800
rect 11878 1724 12014 1734
rect 11772 1452 11854 1462
rect 11528 1440 11610 1450
rect 11610 1374 11772 1408
rect 11772 1362 11854 1372
rect 11528 1350 11610 1360
rect 11654 1278 11736 1288
rect 11914 1278 12014 1724
rect 11890 1268 12014 1278
rect 11736 1214 11890 1248
rect 11654 1188 11736 1198
rect 11972 1188 12014 1268
rect 11890 1178 12014 1188
rect 11914 1174 12014 1178
rect 12606 934 12734 944
rect 11670 922 11794 932
rect 11794 796 12606 906
rect 11670 780 11794 790
rect 12734 796 12744 906
rect 12606 770 12734 780
rect 14260 640 14398 5556
rect 16272 5512 18062 5600
rect 18588 5542 18786 5546
rect 18588 5540 18798 5542
rect 17024 5274 17120 5284
rect 14886 5256 14982 5266
rect 17120 5172 17126 5252
rect 17024 5162 17126 5172
rect 14886 5132 14982 5142
rect 14890 2420 14974 5132
rect 16228 2444 16346 2454
rect 14890 2410 15008 2420
rect 14890 2296 14912 2410
rect 17038 2412 17126 5162
rect 16346 2340 17126 2412
rect 16228 2312 16346 2322
rect 14890 2286 15008 2296
rect 14890 2278 14974 2286
rect 17948 1006 18052 5512
rect 18588 5442 19636 5540
rect 22830 5490 23586 5614
rect 26466 5532 26634 5534
rect 26002 5516 26106 5524
rect 22466 5456 22602 5470
rect 18588 5342 18798 5442
rect 21432 5382 22602 5456
rect 18598 2220 18798 5342
rect 21510 5144 21636 5154
rect 19350 5118 19464 5128
rect 19464 5004 19478 5090
rect 21510 5010 21636 5020
rect 19350 4994 19478 5004
rect 19378 2542 19478 4994
rect 20756 2596 20882 2606
rect 21526 2602 21626 5010
rect 19378 2532 19492 2542
rect 21306 2594 21626 2602
rect 20882 2484 21626 2594
rect 20756 2462 20882 2472
rect 21306 2470 21626 2484
rect 19378 2408 19492 2418
rect 18566 2210 18812 2220
rect 18566 1904 18812 1914
rect 18598 1892 18798 1904
rect 22466 1006 22602 5382
rect 22830 3350 23062 5490
rect 25344 5440 26106 5516
rect 25458 5192 25580 5218
rect 23292 5178 23408 5188
rect 23408 5058 23420 5174
rect 22812 2700 23082 3350
rect 22812 2552 22840 2700
rect 23046 2552 23082 2700
rect 23292 2674 23420 5058
rect 25458 5068 25472 5192
rect 25568 5068 25580 5192
rect 25458 2884 25580 5068
rect 25458 2712 25570 2884
rect 24946 2702 25570 2712
rect 23268 2642 23694 2674
rect 23268 2522 23556 2642
rect 23672 2522 23694 2642
rect 25042 2606 25570 2702
rect 24946 2568 25042 2578
rect 23268 2486 23694 2522
rect 22840 2446 23046 2456
rect 17930 746 22724 1006
rect 21716 672 21944 682
rect 22572 680 22724 746
rect 14260 632 16932 640
rect 14260 596 16988 632
rect 18528 618 18774 628
rect 14260 462 18528 596
rect 14260 456 16426 462
rect 16816 412 18528 462
rect 20880 602 21008 612
rect 18774 458 20880 596
rect 21008 458 21716 596
rect 18774 412 21716 458
rect 18528 312 18774 322
rect 20830 -810 21046 412
rect 21716 330 21944 340
rect 22542 670 22770 680
rect 26002 548 26106 5440
rect 26466 5386 27300 5532
rect 30912 5616 30994 5728
rect 30594 5604 30994 5616
rect 30440 5564 30994 5604
rect 30440 5560 30978 5564
rect 30440 5556 30678 5560
rect 30362 5516 30440 5526
rect 30648 5498 30742 5506
rect 30590 5496 30742 5498
rect 30196 5486 30328 5496
rect 29410 5454 29480 5456
rect 28640 5394 29480 5454
rect 26466 1490 26634 5386
rect 27128 4902 27276 4914
rect 27128 4806 27144 4902
rect 27128 3286 27276 4806
rect 28788 4880 28916 4890
rect 28788 4754 28916 4764
rect 27020 3206 27276 3286
rect 27020 2628 27168 3206
rect 28418 2648 28546 2658
rect 27020 2618 27186 2628
rect 27020 2492 27052 2618
rect 28818 2624 28906 4754
rect 29410 4290 29480 5394
rect 30472 5486 30742 5496
rect 30328 5350 30472 5422
rect 30196 5314 30328 5324
rect 30604 5324 30742 5486
rect 30472 5314 30742 5324
rect 29408 4198 29480 4290
rect 29408 3298 29478 4198
rect 28546 2558 28906 2624
rect 28418 2522 28546 2532
rect 27052 2438 27186 2448
rect 26466 1480 26694 1490
rect 26466 1164 26694 1174
rect 29332 816 29550 3298
rect 30648 3076 30742 5314
rect 30564 3066 30742 3076
rect 30302 3042 30412 3052
rect 30412 2938 30564 3024
rect 30674 2982 30742 3066
rect 30564 2926 30674 2936
rect 30302 2902 30412 2912
rect 30454 2752 30512 2762
rect 30872 2728 30928 2730
rect 30512 2680 30928 2728
rect 30454 2656 30512 2666
rect 29332 548 29542 816
rect 30872 634 30928 2680
rect 22770 406 29542 548
rect 29332 396 29542 406
rect 30862 468 30942 634
rect 22542 328 22770 338
rect 26496 188 26744 198
rect 26496 -20 26744 -10
rect 26544 -810 26682 -20
rect 20830 -822 26712 -810
rect 30862 -822 30936 468
rect 20830 -1030 30936 -822
rect 20830 -1056 26712 -1030
rect 20830 -1060 21046 -1056
<< via2 >>
rect 11632 6068 11722 6090
rect 11632 6002 11642 6068
rect 11642 6002 11696 6068
rect 11696 6002 11722 6068
rect 11632 5972 11722 6002
rect 11880 6076 11970 6092
rect 11880 5986 11900 6076
rect 11900 5986 11962 6076
rect 11962 5986 11970 6076
rect 11620 5752 11710 5774
rect 11880 5974 11970 5986
rect 11620 5686 11640 5752
rect 11640 5686 11694 5752
rect 11694 5686 11710 5752
rect 11620 5656 11710 5686
rect 11882 5758 11972 5778
rect 11882 5668 11902 5758
rect 11902 5668 11964 5758
rect 11964 5668 11972 5758
rect 11626 5428 11716 5458
rect 11882 5660 11972 5668
rect 11626 5362 11650 5428
rect 11650 5362 11704 5428
rect 11704 5362 11716 5428
rect 11626 5340 11716 5362
rect 11880 5438 11970 5458
rect 11880 5348 11894 5438
rect 11894 5348 11956 5438
rect 11956 5348 11970 5438
rect 11880 5340 11970 5348
rect 11638 5106 11728 5132
rect 11638 5040 11646 5106
rect 11646 5040 11700 5106
rect 11700 5040 11728 5106
rect 11638 5014 11728 5040
rect 11876 5116 11966 5132
rect 11876 5026 11888 5116
rect 11888 5026 11950 5116
rect 11950 5026 11966 5116
rect 11876 5014 11966 5026
rect 11626 4786 11716 4816
rect 11626 4720 11650 4786
rect 11650 4720 11704 4786
rect 11704 4720 11716 4786
rect 11626 4698 11716 4720
rect 11880 4800 11970 4812
rect 11880 4710 11892 4800
rect 11892 4710 11954 4800
rect 11954 4710 11970 4800
rect 11880 4694 11970 4710
rect 11628 4464 11714 4488
rect 11628 4398 11646 4464
rect 11646 4398 11700 4464
rect 11700 4398 11714 4464
rect 11628 4374 11714 4398
rect 11876 4476 11962 4490
rect 11876 4386 11888 4476
rect 11888 4386 11950 4476
rect 11950 4386 11962 4476
rect 11876 4376 11962 4386
rect 11628 4140 11726 4164
rect 11628 4080 11638 4140
rect 11638 4080 11694 4140
rect 11694 4080 11726 4140
rect 11628 4066 11726 4080
rect 11870 4148 11966 4166
rect 11870 4078 11890 4148
rect 11890 4078 11944 4148
rect 11944 4078 11966 4148
rect 11870 4068 11966 4078
rect 11630 3828 11720 3856
rect 11874 3840 11964 3860
rect 11630 3762 11642 3828
rect 11642 3762 11696 3828
rect 11696 3762 11720 3828
rect 11630 3738 11720 3762
rect 11874 3750 11896 3840
rect 11896 3750 11958 3840
rect 11958 3750 11964 3840
rect 11874 3742 11964 3750
rect 11626 3512 11716 3534
rect 11626 3446 11642 3512
rect 11642 3446 11696 3512
rect 11696 3446 11716 3512
rect 11626 3416 11716 3446
rect 11872 3522 11962 3532
rect 11872 3432 11888 3522
rect 11888 3432 11950 3522
rect 11950 3432 11962 3522
rect 11618 3186 11708 3214
rect 11872 3414 11962 3432
rect 11618 3120 11638 3186
rect 11638 3120 11692 3186
rect 11692 3120 11708 3186
rect 11618 3096 11708 3120
rect 11880 3200 11970 3212
rect 11880 3110 11894 3200
rect 11894 3110 11956 3200
rect 11956 3110 11970 3200
rect 11880 3094 11970 3110
<< metal3 >>
rect 11622 6090 11732 6095
rect 11622 5972 11632 6090
rect 11722 6078 11732 6090
rect 11870 6092 11980 6097
rect 11870 6078 11880 6092
rect 11722 5988 11880 6078
rect 11722 5972 11732 5988
rect 11622 5967 11732 5972
rect 11870 5974 11880 5988
rect 11970 5974 11980 6092
rect 11870 5969 11980 5974
rect 11610 5774 11720 5779
rect 11610 5656 11620 5774
rect 11710 5762 11720 5774
rect 11872 5778 11982 5783
rect 11872 5762 11882 5778
rect 11710 5672 11882 5762
rect 11710 5656 11720 5672
rect 11610 5651 11720 5656
rect 11872 5660 11882 5672
rect 11972 5660 11982 5778
rect 11872 5655 11982 5660
rect 11616 5458 11726 5463
rect 11616 5340 11626 5458
rect 11716 5440 11726 5458
rect 11870 5458 11980 5463
rect 11870 5440 11880 5458
rect 11716 5350 11880 5440
rect 11716 5340 11726 5350
rect 11616 5335 11726 5340
rect 11870 5340 11880 5350
rect 11970 5340 11980 5458
rect 11870 5335 11980 5340
rect 11628 5132 11738 5137
rect 11628 5014 11638 5132
rect 11728 5122 11738 5132
rect 11866 5132 11976 5137
rect 11866 5122 11876 5132
rect 11728 5032 11876 5122
rect 11728 5014 11738 5032
rect 11628 5009 11738 5014
rect 11866 5014 11876 5032
rect 11966 5014 11976 5132
rect 11866 5009 11976 5014
rect 11616 4816 11726 4821
rect 11616 4698 11626 4816
rect 11716 4786 11726 4816
rect 11870 4812 11980 4817
rect 11870 4786 11880 4812
rect 11716 4718 11880 4786
rect 11716 4698 11726 4718
rect 11616 4693 11726 4698
rect 11870 4694 11880 4718
rect 11970 4694 11980 4812
rect 11870 4689 11980 4694
rect 11618 4488 11724 4493
rect 11618 4374 11628 4488
rect 11714 4464 11724 4488
rect 11866 4490 11972 4495
rect 11866 4464 11876 4490
rect 11714 4400 11876 4464
rect 11714 4374 11724 4400
rect 11618 4369 11724 4374
rect 11866 4376 11876 4400
rect 11962 4376 11972 4490
rect 11866 4371 11972 4376
rect 11618 4164 11736 4169
rect 11618 4066 11628 4164
rect 11726 4156 11736 4164
rect 11860 4166 11976 4171
rect 11860 4156 11870 4166
rect 11726 4078 11870 4156
rect 11726 4066 11736 4078
rect 11618 4061 11736 4066
rect 11860 4068 11870 4078
rect 11966 4068 11976 4166
rect 11860 4063 11976 4068
rect 11620 3856 11730 3861
rect 11620 3738 11630 3856
rect 11720 3830 11730 3856
rect 11864 3860 11974 3865
rect 11864 3830 11874 3860
rect 11720 3766 11874 3830
rect 11720 3738 11730 3766
rect 11620 3733 11730 3738
rect 11864 3742 11874 3766
rect 11964 3742 11974 3860
rect 11864 3737 11974 3742
rect 11616 3534 11726 3539
rect 11616 3416 11626 3534
rect 11716 3508 11726 3534
rect 11862 3532 11972 3537
rect 11862 3508 11872 3532
rect 11716 3444 11872 3508
rect 11716 3416 11726 3444
rect 11616 3411 11726 3416
rect 11862 3414 11872 3444
rect 11962 3414 11972 3532
rect 11862 3409 11972 3414
rect 11608 3214 11718 3219
rect 11608 3096 11618 3214
rect 11708 3200 11718 3214
rect 11870 3212 11980 3217
rect 11870 3200 11880 3212
rect 11708 3138 11880 3200
rect 11708 3096 11718 3138
rect 11608 3091 11718 3096
rect 11870 3094 11880 3138
rect 11970 3094 11980 3212
rect 11870 3089 11980 3094
use sky130_fd_pr__res_generic_po_4WEV9M  R1
timestamp 1754378775
transform 1 0 22662 0 1 103
box -266 -761 266 761
use sky130_fd_pr__res_generic_po_4WEV9M  R4
timestamp 1754378775
transform 1 0 21844 0 1 127
box -266 -761 266 761
use inv_layout_tt  x1
timestamp 1755205548
transform 1 0 15908 0 1 3430
box -1072 -1780 500 -190
use inv_layout_tt  x2
timestamp 1755205548
transform 1 0 20414 0 1 3586
box -1072 -1780 500 -190
use inv_layout_tt  x3
timestamp 1755205548
transform 1 0 24602 0 1 3684
box -1072 -1780 500 -190
use dac_inside_tt_v2  x4
timestamp 1755204415
transform 1 0 18440 0 1 5778
box 204 -1268 3482 1496
use inv_layout_tt  x5
timestamp 1755205548
transform 1 0 28088 0 1 3618
box -1072 -1780 500 -190
use dac_inside_tt_v2  x6
timestamp 1755204415
transform 1 0 22396 0 1 5844
box 204 -1268 3482 1496
use dac_inside_tt  x8
timestamp 1755120335
transform 1 0 26466 0 1 6230
box 484 -1844 2714 456
use dac_inside_tt_v2  x9
timestamp 1755204415
transform 1 0 13956 0 1 5914
box 204 -1268 3482 1496
use sky130_fd_pr__pfet_01v8_4YM9M3  XM4
timestamp 1754378775
transform 1 0 11734 0 1 4593
box -344 -1701 344 1701
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM15
timestamp 1754378775
transform 1 0 30397 0 1 5379
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM18
timestamp 1754378775
transform 1 0 30487 0 1 2831
box -285 -469 285 469
use sky130_fd_pr__nfet_01v8_93A3ZJ  XM31
timestamp 1754378775
transform 1 0 11746 0 1 1585
box -344 -653 344 653
<< labels >>
flabel metal1 11818 7586 12018 7786 0 FreeSans 256 0 0 0 Vdd
port 0 nsew
flabel metal1 11902 576 12102 776 0 FreeSans 256 0 0 0 Vss
port 1 nsew
flabel metal1 20854 438 21054 638 0 FreeSans 256 0 0 0 Vout1
port 6 nsew
flabel metal1 23088 414 23288 614 0 FreeSans 256 0 0 0 Vout2
port 7 nsew
flabel metal1 14492 2246 14692 2446 0 FreeSans 256 0 0 0 Vin4
port 5 nsew
flabel metal1 19024 2398 19224 2598 0 FreeSans 256 0 0 0 Vin3
port 4 nsew
flabel metal1 23280 1994 23480 2194 0 FreeSans 256 0 0 0 Vin2
port 3 nsew
flabel metal1 26782 2022 26982 2222 0 FreeSans 256 0 0 0 Vin1
port 2 nsew
rlabel metal2 30674 3912 30710 4012 1 net33
rlabel metal1 13584 6474 13712 6618 1 Vg
<< end >>
