
* expanding   symbol:  /home/eserlis/one_class_tt_official.sym # of pins=10
** sym_path: /home/eserlis/one_class_tt_official.sym
** sch_path: /home/eserlis/one_class_tt_official.sch
.subckt one_class_tt_official Vdd Vss Vr Vin4 Vin3 Vin2 Vin1 En Iout0 Iout1
*.iopin Vdd
*.iopin Vr
*.iopin Vss
*.iopin Vin3
*.iopin Vin2
*.iopin Vin1
*.iopin Vin4
*.iopin En
*.iopin Iout0
*.iopin Iout1
x5 Vdd Iout00 Vr Vdac0 Ibias Vss bump_final_tt
x2 Vdd Iout01 Vr Vdac0 Iout00 Vss bump_final_tt
x6 Vdd Iout10 Vref4 Vdac1 Ibias Vss bump_final_tt
x7 Vdd Iout11 Vref4 Vdac1 Iout10 Vss bump_final_tt
x11 Vdd En Ibias Vss ref_gen_tt
x3 Vref2 Vdd Vref1 Vss Vref3 Vref4 vol_ref_gen_tt
x1 Vdd Vss Vin1dac Vin2dac Vin3dac Vin4dac Vdac0 Vdac1 dac_tt
x4 Iout11 Iclass1 Vss ccm_nmos_tt
x8 Iout01 Iclass0 Vss ccm_nmos_tt
x12 Vdd Vss Iout0 Iout1 Iclass0 Iclass1 Ibias wta_pmos_tt
x9 Vss Vdd Vin3dac Vin3 inv_layout_tt
x10 Vss Vdd Vin4dac Vin4 inv_layout_tt
x13 Vss Vdd Vin1dac Vin1 inv_layout_tt
x14 Vss Vdd Vin2dac Vin2 inv_layout_tt
R964 Vdd.n409 Vdd.n406 6783.53
R965 Vdd.n412 Vdd.n405 6783.53
R966 Vdd.n60 Vdd.n59 2975.29
R967 Vdd.n62 Vdd.n53 2975.29
R968 Vdd.n31 Vdd.n30 2975.29
R969 Vdd.n83 Vdd.n29 2975.29
R970 Vdd.n17 Vdd.n16 2505.88
R971 Vdd.n19 Vdd.n13 2505.88
R972 Vdd.n373 Vdd.n371 2227.06
R973 Vdd.n376 Vdd.n375 2227.06
R974 Vdd.n358 Vdd.n356 2227.06
R975 Vdd.n365 Vdd.n354 2227.06
R976 Vdd.n321 Vdd.n310 2227.06
R977 Vdd.n314 Vdd.n312 2227.06
R978 Vdd.n332 Vdd.n331 2227.06
R979 Vdd.n329 Vdd.n327 2227.06
R980 Vdd.n225 Vdd.n219 2227.06
R981 Vdd.n222 Vdd.n220 2227.06
R982 Vdd.n214 Vdd.n208 2227.06
R983 Vdd.n211 Vdd.n209 2227.06
R984 Vdd.n202 Vdd.n199 2227.06
R985 Vdd.n253 Vdd.n197 2227.06
R986 Vdd.n235 Vdd.n234 2227.06
R987 Vdd.n237 Vdd.n231 2227.06
R988 Vdd.n275 Vdd.n264 2227.06
R989 Vdd.n268 Vdd.n266 2227.06
R990 Vdd.n286 Vdd.n285 2227.06
R991 Vdd.n283 Vdd.n281 2227.06
R992 Vdd.n136 Vdd.n135 1912.94
R993 Vdd.n138 Vdd.n132 1912.94
R994 Vdd.n150 Vdd.n149 1912.94
R995 Vdd.n152 Vdd.n146 1912.94
R996 Vdd.n176 Vdd.n175 1912.94
R997 Vdd.n178 Vdd.n172 1912.94
R998 Vdd.n188 Vdd.n187 1912.94
R999 Vdd.n190 Vdd.n184 1912.94
R1000 Vdd.n163 Vdd.n162 1912.94
R1001 Vdd.n165 Vdd.n159 1912.94
R1002 Vdd.n123 Vdd.n122 1912.94
R1003 Vdd.n125 Vdd.n119 1912.94
R1004 Vdd.n94 Vdd.n93 1912.94
R1005 Vdd.n96 Vdd.n90 1912.94
R1006 Vdd.n108 Vdd.n107 1912.94
R1007 Vdd.n110 Vdd.n104 1912.94
R1008 Vdd.n687 Vdd.n671 1807.06
R1009 Vdd.n680 Vdd.n676 1807.06
R1010 Vdd.n611 Vdd.n595 1807.06
R1011 Vdd.n604 Vdd.n600 1807.06
R1012 Vdd.n535 Vdd.n519 1807.06
R1013 Vdd.n528 Vdd.n524 1807.06
R1014 Vdd.n460 Vdd.n444 1807.06
R1015 Vdd.n453 Vdd.n449 1807.06
R1016 Vdd.n739 Vdd.n738 1771.76
R1017 Vdd.n751 Vdd.n750 1771.76
R1018 Vdd.n736 Vdd.n731 1771.76
R1019 Vdd.n748 Vdd.n743 1771.76
R1020 Vdd.n657 Vdd.n653 1771.76
R1021 Vdd.n664 Vdd.n648 1771.76
R1022 Vdd.n711 Vdd.n695 1771.76
R1023 Vdd.n704 Vdd.n700 1771.76
R1024 Vdd.n635 Vdd.n619 1771.76
R1025 Vdd.n628 Vdd.n624 1771.76
R1026 Vdd.n581 Vdd.n577 1771.76
R1027 Vdd.n588 Vdd.n572 1771.76
R1028 Vdd.n505 Vdd.n501 1771.76
R1029 Vdd.n512 Vdd.n496 1771.76
R1030 Vdd.n559 Vdd.n543 1771.76
R1031 Vdd.n552 Vdd.n548 1771.76
R1032 Vdd.n430 Vdd.n426 1771.76
R1033 Vdd.n437 Vdd.n421 1771.76
R1034 Vdd.n484 Vdd.n468 1771.76
R1035 Vdd.n477 Vdd.n473 1771.76
R1036 Vdd.n59 Vdd.n55 1736.47
R1037 Vdd.n55 Vdd.n53 1736.47
R1038 Vdd.n68 Vdd.n44 1736.47
R1039 Vdd.n68 Vdd.n67 1736.47
R1040 Vdd.n67 Vdd.n66 1736.47
R1041 Vdd.n66 Vdd.n37 1736.47
R1042 Vdd.n30 Vdd.n28 1736.47
R1043 Vdd.n83 Vdd.n28 1736.47
R1044 Vdd.n43 Vdd.n42 1736.47
R1045 Vdd.n42 Vdd.n33 1736.47
R1046 Vdd.n76 Vdd.n33 1736.47
R1047 Vdd.n76 Vdd.n75 1736.47
R1048 Vdd.n410 Vdd.n405 1720.44
R1049 Vdd.n411 Vdd.n406 1720.44
R1050 Vdd.n371 Vdd.n350 1408.24
R1051 Vdd.n369 Vdd.n351 1408.24
R1052 Vdd.n370 Vdd.n369 1408.24
R1053 Vdd.n360 Vdd.n359 1408.24
R1054 Vdd.n360 Vdd.n351 1408.24
R1055 Vdd.n366 Vdd.n365 1408.24
R1056 Vdd.n376 Vdd.n366 1408.24
R1057 Vdd.n356 Vdd.n350 1408.24
R1058 Vdd.n322 Vdd.n321 1408.24
R1059 Vdd.n312 Vdd.n306 1408.24
R1060 Vdd.n316 Vdd.n315 1408.24
R1061 Vdd.n316 Vdd.n307 1408.24
R1062 Vdd.n325 Vdd.n307 1408.24
R1063 Vdd.n326 Vdd.n325 1408.24
R1064 Vdd.n332 Vdd.n322 1408.24
R1065 Vdd.n327 Vdd.n306 1408.24
R1066 Vdd.n249 Vdd.n200 1408.24
R1067 Vdd.n250 Vdd.n249 1408.24
R1068 Vdd.n276 Vdd.n275 1408.24
R1069 Vdd.n266 Vdd.n260 1408.24
R1070 Vdd.n270 Vdd.n269 1408.24
R1071 Vdd.n270 Vdd.n261 1408.24
R1072 Vdd.n279 Vdd.n261 1408.24
R1073 Vdd.n280 Vdd.n279 1408.24
R1074 Vdd.n286 Vdd.n276 1408.24
R1075 Vdd.n281 Vdd.n260 1408.24
R1076 Vdd.n5 Vdd.n3 1383.53
R1077 Vdd.n8 Vdd.n2 1383.53
R1078 Vdd.n72 Vdd.n43 1238.82
R1079 Vdd.n72 Vdd.n44 1238.82
R1080 Vdd.n60 Vdd.n44 1238.82
R1081 Vdd.n62 Vdd.n37 1238.82
R1082 Vdd.n40 Vdd.n33 1238.82
R1083 Vdd.n67 Vdd.n40 1238.82
R1084 Vdd.n67 Vdd.n50 1238.82
R1085 Vdd.n55 Vdd.n50 1238.82
R1086 Vdd.n80 Vdd.n28 1238.82
R1087 Vdd.n80 Vdd.n33 1238.82
R1088 Vdd.n75 Vdd.n29 1238.82
R1089 Vdd.n75 Vdd.n74 1238.82
R1090 Vdd.n74 Vdd.n37 1238.82
R1091 Vdd.n43 Vdd.n31 1238.82
R1092 Vdd.n739 Vdd.n728 1069.41
R1093 Vdd.n751 Vdd.n728 1069.41
R1094 Vdd.n731 Vdd.n724 1069.41
R1095 Vdd.n743 Vdd.n724 1069.41
R1096 Vdd.n732 Vdd.n730 1069.41
R1097 Vdd.n732 Vdd.n725 1069.41
R1098 Vdd.n744 Vdd.n725 1069.41
R1099 Vdd.n744 Vdd.n742 1069.41
R1100 Vdd.n654 Vdd.n647 1069.41
R1101 Vdd.n664 Vdd.n647 1069.41
R1102 Vdd.n657 Vdd.n651 1069.41
R1103 Vdd.n661 Vdd.n651 1069.41
R1104 Vdd.n680 Vdd.n674 1069.41
R1105 Vdd.n684 Vdd.n674 1069.41
R1106 Vdd.n677 Vdd.n670 1069.41
R1107 Vdd.n687 Vdd.n670 1069.41
R1108 Vdd.n704 Vdd.n698 1069.41
R1109 Vdd.n708 Vdd.n698 1069.41
R1110 Vdd.n701 Vdd.n694 1069.41
R1111 Vdd.n711 Vdd.n694 1069.41
R1112 Vdd.n628 Vdd.n622 1069.41
R1113 Vdd.n632 Vdd.n622 1069.41
R1114 Vdd.n625 Vdd.n618 1069.41
R1115 Vdd.n635 Vdd.n618 1069.41
R1116 Vdd.n578 Vdd.n571 1069.41
R1117 Vdd.n588 Vdd.n571 1069.41
R1118 Vdd.n581 Vdd.n575 1069.41
R1119 Vdd.n585 Vdd.n575 1069.41
R1120 Vdd.n604 Vdd.n598 1069.41
R1121 Vdd.n608 Vdd.n598 1069.41
R1122 Vdd.n601 Vdd.n594 1069.41
R1123 Vdd.n611 Vdd.n594 1069.41
R1124 Vdd.n502 Vdd.n495 1069.41
R1125 Vdd.n512 Vdd.n495 1069.41
R1126 Vdd.n505 Vdd.n499 1069.41
R1127 Vdd.n509 Vdd.n499 1069.41
R1128 Vdd.n528 Vdd.n522 1069.41
R1129 Vdd.n532 Vdd.n522 1069.41
R1130 Vdd.n525 Vdd.n518 1069.41
R1131 Vdd.n535 Vdd.n518 1069.41
R1132 Vdd.n552 Vdd.n546 1069.41
R1133 Vdd.n556 Vdd.n546 1069.41
R1134 Vdd.n549 Vdd.n542 1069.41
R1135 Vdd.n559 Vdd.n542 1069.41
R1136 Vdd.n427 Vdd.n420 1069.41
R1137 Vdd.n437 Vdd.n420 1069.41
R1138 Vdd.n430 Vdd.n424 1069.41
R1139 Vdd.n434 Vdd.n424 1069.41
R1140 Vdd.n453 Vdd.n447 1069.41
R1141 Vdd.n457 Vdd.n447 1069.41
R1142 Vdd.n450 Vdd.n443 1069.41
R1143 Vdd.n460 Vdd.n443 1069.41
R1144 Vdd.n477 Vdd.n471 1069.41
R1145 Vdd.n481 Vdd.n471 1069.41
R1146 Vdd.n474 Vdd.n467 1069.41
R1147 Vdd.n484 Vdd.n467 1069.41
R1148 Vdd.n373 Vdd.n370 818.823
R1149 Vdd.n375 Vdd.n370 818.823
R1150 Vdd.n359 Vdd.n358 818.823
R1151 Vdd.n359 Vdd.n354 818.823
R1152 Vdd.n382 Vdd.n350 818.823
R1153 Vdd.n382 Vdd.n351 818.823
R1154 Vdd.n380 Vdd.n351 818.823
R1155 Vdd.n380 Vdd.n366 818.823
R1156 Vdd.n315 Vdd.n314 818.823
R1157 Vdd.n315 Vdd.n310 818.823
R1158 Vdd.n338 Vdd.n306 818.823
R1159 Vdd.n338 Vdd.n307 818.823
R1160 Vdd.n336 Vdd.n307 818.823
R1161 Vdd.n336 Vdd.n322 818.823
R1162 Vdd.n329 Vdd.n326 818.823
R1163 Vdd.n331 Vdd.n326 818.823
R1164 Vdd.n245 Vdd.n200 818.823
R1165 Vdd.n200 Vdd.n197 818.823
R1166 Vdd.n250 Vdd.n199 818.823
R1167 Vdd.n251 Vdd.n250 818.823
R1168 Vdd.n269 Vdd.n268 818.823
R1169 Vdd.n269 Vdd.n264 818.823
R1170 Vdd.n292 Vdd.n260 818.823
R1171 Vdd.n292 Vdd.n261 818.823
R1172 Vdd.n290 Vdd.n261 818.823
R1173 Vdd.n290 Vdd.n276 818.823
R1174 Vdd.n283 Vdd.n280 818.823
R1175 Vdd.n285 Vdd.n280 818.823
R1176 Vdd.n673 Vdd.n670 737.648
R1177 Vdd.n674 Vdd.n673 737.648
R1178 Vdd.n597 Vdd.n594 737.648
R1179 Vdd.n598 Vdd.n597 737.648
R1180 Vdd.n521 Vdd.n518 737.648
R1181 Vdd.n522 Vdd.n521 737.648
R1182 Vdd.n446 Vdd.n443 737.648
R1183 Vdd.n447 Vdd.n446 737.648
R1184 Vdd.n408 Vdd.n407 723.577
R1185 Vdd.n408 Vdd.n404 723.577
R1186 Vdd.n413 Vdd.n404 723.577
R1187 Vdd.n407 Vdd.n403 717.177
R1188 Vdd.n755 Vdd.n725 702.354
R1189 Vdd.n755 Vdd.n728 702.354
R1190 Vdd.n738 Vdd.n730 702.354
R1191 Vdd.n757 Vdd.n724 702.354
R1192 Vdd.n757 Vdd.n725 702.354
R1193 Vdd.n736 Vdd.n730 702.354
R1194 Vdd.n748 Vdd.n742 702.354
R1195 Vdd.n750 Vdd.n742 702.354
R1196 Vdd.n650 Vdd.n647 702.354
R1197 Vdd.n651 Vdd.n650 702.354
R1198 Vdd.n697 Vdd.n694 702.354
R1199 Vdd.n698 Vdd.n697 702.354
R1200 Vdd.n621 Vdd.n618 702.354
R1201 Vdd.n622 Vdd.n621 702.354
R1202 Vdd.n574 Vdd.n571 702.354
R1203 Vdd.n575 Vdd.n574 702.354
R1204 Vdd.n498 Vdd.n495 702.354
R1205 Vdd.n499 Vdd.n498 702.354
R1206 Vdd.n545 Vdd.n542 702.354
R1207 Vdd.n546 Vdd.n545 702.354
R1208 Vdd.n423 Vdd.n420 702.354
R1209 Vdd.n424 Vdd.n423 702.354
R1210 Vdd.n470 Vdd.n467 702.354
R1211 Vdd.n471 Vdd.n470 702.354
R1212 Vdd.n19 Vdd.n18 611.4
R1213 Vdd.n16 Vdd.n14 611.4
R1214 Vdd.n223 Vdd.n219 546.558
R1215 Vdd.n224 Vdd.n220 546.558
R1216 Vdd.n212 Vdd.n208 546.558
R1217 Vdd.n213 Vdd.n209 546.558
R1218 Vdd.n237 Vdd.n236 546.558
R1219 Vdd.n234 Vdd.n232 546.558
R1220 Vdd.n135 Vdd.n133 543.497
R1221 Vdd.n138 Vdd.n137 543.497
R1222 Vdd.n149 Vdd.n147 543.497
R1223 Vdd.n152 Vdd.n151 543.497
R1224 Vdd.n175 Vdd.n173 543.497
R1225 Vdd.n178 Vdd.n177 543.497
R1226 Vdd.n187 Vdd.n185 543.497
R1227 Vdd.n190 Vdd.n189 543.497
R1228 Vdd.n162 Vdd.n160 543.497
R1229 Vdd.n165 Vdd.n164 543.497
R1230 Vdd.n122 Vdd.n120 543.497
R1231 Vdd.n125 Vdd.n124 543.497
R1232 Vdd.n93 Vdd.n91 543.497
R1233 Vdd.n96 Vdd.n95 543.497
R1234 Vdd.n107 Vdd.n105 543.497
R1235 Vdd.n110 Vdd.n109 543.497
R1236 Vdd.n656 Vdd.n649 535.038
R1237 Vdd.n663 Vdd.n649 535.038
R1238 Vdd.n703 Vdd.n696 535.038
R1239 Vdd.n710 Vdd.n696 535.038
R1240 Vdd.n627 Vdd.n620 535.038
R1241 Vdd.n634 Vdd.n620 535.038
R1242 Vdd.n580 Vdd.n573 535.038
R1243 Vdd.n587 Vdd.n573 535.038
R1244 Vdd.n504 Vdd.n497 535.038
R1245 Vdd.n511 Vdd.n497 535.038
R1246 Vdd.n551 Vdd.n544 535.038
R1247 Vdd.n558 Vdd.n544 535.038
R1248 Vdd.n429 Vdd.n422 535.038
R1249 Vdd.n436 Vdd.n422 535.038
R1250 Vdd.n476 Vdd.n469 535.038
R1251 Vdd.n483 Vdd.n469 535.038
R1252 Vdd.n679 Vdd.n672 515.861
R1253 Vdd.n686 Vdd.n672 515.861
R1254 Vdd.n603 Vdd.n596 515.861
R1255 Vdd.n610 Vdd.n596 515.861
R1256 Vdd.n527 Vdd.n520 515.861
R1257 Vdd.n534 Vdd.n520 515.861
R1258 Vdd.n452 Vdd.n445 515.861
R1259 Vdd.n459 Vdd.n445 515.861
R1260 Vdd.n655 Vdd.n653 432.829
R1261 Vdd.n662 Vdd.n648 432.829
R1262 Vdd.n702 Vdd.n700 432.829
R1263 Vdd.n709 Vdd.n695 432.829
R1264 Vdd.n626 Vdd.n624 432.829
R1265 Vdd.n633 Vdd.n619 432.829
R1266 Vdd.n579 Vdd.n577 432.829
R1267 Vdd.n586 Vdd.n572 432.829
R1268 Vdd.n503 Vdd.n501 432.829
R1269 Vdd.n510 Vdd.n496 432.829
R1270 Vdd.n550 Vdd.n548 432.829
R1271 Vdd.n557 Vdd.n543 432.829
R1272 Vdd.n428 Vdd.n426 432.829
R1273 Vdd.n435 Vdd.n421 432.829
R1274 Vdd.n475 Vdd.n473 432.829
R1275 Vdd.n482 Vdd.n468 432.829
R1276 Vdd.n678 Vdd.n676 424.014
R1277 Vdd.n685 Vdd.n671 424.014
R1278 Vdd.n602 Vdd.n600 424.014
R1279 Vdd.n609 Vdd.n595 424.014
R1280 Vdd.n526 Vdd.n524 424.014
R1281 Vdd.n533 Vdd.n519 424.014
R1282 Vdd.n451 Vdd.n449 424.014
R1283 Vdd.n458 Vdd.n444 424.014
R1284 Vdd.n357 Vdd.n352 382.205
R1285 Vdd.n381 Vdd.n352 382.205
R1286 Vdd.n381 Vdd.n353 382.205
R1287 Vdd.n374 Vdd.n353 382.205
R1288 Vdd.n313 Vdd.n308 382.205
R1289 Vdd.n337 Vdd.n308 382.205
R1290 Vdd.n337 Vdd.n309 382.205
R1291 Vdd.n330 Vdd.n309 382.205
R1292 Vdd.n267 Vdd.n262 382.205
R1293 Vdd.n291 Vdd.n262 382.205
R1294 Vdd.n291 Vdd.n263 382.205
R1295 Vdd.n284 Vdd.n263 382.205
R1296 Vdd.n6 Vdd.n2 347.05
R1297 Vdd.n7 Vdd.n3 347.05
R1298 Vdd.n394 Vdd.t0 337.618
R1299 Vdd.n398 Vdd.t4 337.615
R1300 Vdd.t2 Vdd.n396 337.586
R1301 Vdd.t3 Vdd.n395 337.231
R1302 Vdd.n396 Vdd.t3 337.231
R1303 Vdd.n397 Vdd.t2 337.231
R1304 Vdd.t1 Vdd.n392 337.231
R1305 Vdd.n393 Vdd.t1 337.231
R1306 Vdd.t4 Vdd.n397 337.231
R1307 Vdd.t5 Vdd.n394 337.231
R1308 Vdd.n395 Vdd.t5 337.231
R1309 Vdd.t0 Vdd.n393 337.231
R1310 Vdd.n84 Vdd.n27 317.365
R1311 Vdd.n58 Vdd.n48 317.365
R1312 Vdd.n63 Vdd.n52 317.365
R1313 Vdd.n46 Vdd.n45 316.714
R1314 Vdd.n737 Vdd.n726 296.753
R1315 Vdd.n756 Vdd.n726 296.753
R1316 Vdd.n756 Vdd.n727 296.753
R1317 Vdd.n749 Vdd.n727 296.753
R1318 Vdd.n20 Vdd.n12 267.295
R1319 Vdd.n15 Vdd.n12 267.295
R1320 Vdd.n15 Vdd.n11 267.295
R1321 Vdd.n372 Vdd.n348 237.554
R1322 Vdd.n377 Vdd.n367 237.554
R1323 Vdd.n364 Vdd.n363 237.554
R1324 Vdd.n333 Vdd.n323 237.554
R1325 Vdd.n320 Vdd.n319 237.554
R1326 Vdd.n328 Vdd.n304 237.554
R1327 Vdd.n221 Vdd.n217 237.554
R1328 Vdd.n221 Vdd.n218 237.554
R1329 Vdd.n226 Vdd.n218 237.554
R1330 Vdd.n210 Vdd.n206 237.554
R1331 Vdd.n210 Vdd.n207 237.554
R1332 Vdd.n215 Vdd.n207 237.554
R1333 Vdd.n254 Vdd.n196 237.554
R1334 Vdd.n205 Vdd.n204 237.554
R1335 Vdd.n238 Vdd.n230 237.554
R1336 Vdd.n233 Vdd.n230 237.554
R1337 Vdd.n233 Vdd.n229 237.554
R1338 Vdd.n287 Vdd.n277 237.554
R1339 Vdd.n274 Vdd.n273 237.554
R1340 Vdd.n282 Vdd.n258 237.554
R1341 Vdd.n265 Vdd.n257 237.554
R1342 Vdd.n311 Vdd.n303 237.554
R1343 Vdd.n355 Vdd.n347 237.554
R1344 Vdd.n248 Vdd.n247 234.969
R1345 Vdd.n248 Vdd.n198 234.969
R1346 Vdd.n239 Vdd.n229 226.403
R1347 Vdd.n253 Vdd.n252 224.225
R1348 Vdd.n246 Vdd.n202 224.225
R1349 Vdd.n134 Vdd.n131 204.048
R1350 Vdd.n139 Vdd.n131 204.048
R1351 Vdd.n148 Vdd.n145 204.048
R1352 Vdd.n153 Vdd.n145 204.048
R1353 Vdd.n174 Vdd.n171 204.048
R1354 Vdd.n179 Vdd.n171 204.048
R1355 Vdd.n186 Vdd.n183 204.048
R1356 Vdd.n191 Vdd.n183 204.048
R1357 Vdd.n161 Vdd.n158 204.048
R1358 Vdd.n166 Vdd.n158 204.048
R1359 Vdd.n121 Vdd.n118 204.048
R1360 Vdd.n126 Vdd.n118 204.048
R1361 Vdd.n92 Vdd.n89 204.048
R1362 Vdd.n97 Vdd.n89 204.048
R1363 Vdd.n106 Vdd.n103 204.048
R1364 Vdd.n111 Vdd.n103 204.048
R1365 Vdd.n134 Vdd.n130 203.719
R1366 Vdd.n148 Vdd.n144 203.719
R1367 Vdd.n174 Vdd.n170 203.719
R1368 Vdd.n186 Vdd.n182 203.719
R1369 Vdd.n161 Vdd.n157 203.719
R1370 Vdd.n121 Vdd.n117 203.719
R1371 Vdd.n92 Vdd.n88 203.719
R1372 Vdd.n106 Vdd.n102 203.719
R1373 Vdd.n21 Vdd.n11 200.689
R1374 Vdd.n675 Vdd.n667 192.754
R1375 Vdd.n681 Vdd.n675 192.754
R1376 Vdd.n688 Vdd.n669 192.754
R1377 Vdd.n683 Vdd.n669 192.754
R1378 Vdd.n599 Vdd.n591 192.754
R1379 Vdd.n605 Vdd.n599 192.754
R1380 Vdd.n612 Vdd.n593 192.754
R1381 Vdd.n607 Vdd.n593 192.754
R1382 Vdd.n523 Vdd.n515 192.754
R1383 Vdd.n529 Vdd.n523 192.754
R1384 Vdd.n536 Vdd.n517 192.754
R1385 Vdd.n531 Vdd.n517 192.754
R1386 Vdd.n448 Vdd.n440 192.754
R1387 Vdd.n454 Vdd.n448 192.754
R1388 Vdd.n461 Vdd.n442 192.754
R1389 Vdd.n456 Vdd.n442 192.754
R1390 Vdd.n740 Vdd.n729 188.988
R1391 Vdd.n752 Vdd.n741 188.988
R1392 Vdd.n747 Vdd.n722 188.988
R1393 Vdd.n735 Vdd.n721 188.988
R1394 Vdd.n665 Vdd.n646 188.988
R1395 Vdd.n660 Vdd.n646 188.988
R1396 Vdd.n658 Vdd.n652 188.988
R1397 Vdd.n652 Vdd.n645 188.988
R1398 Vdd.n699 Vdd.n691 188.988
R1399 Vdd.n705 Vdd.n699 188.988
R1400 Vdd.n712 Vdd.n693 188.988
R1401 Vdd.n707 Vdd.n693 188.988
R1402 Vdd.n623 Vdd.n615 188.988
R1403 Vdd.n629 Vdd.n623 188.988
R1404 Vdd.n636 Vdd.n617 188.988
R1405 Vdd.n631 Vdd.n617 188.988
R1406 Vdd.n589 Vdd.n570 188.988
R1407 Vdd.n584 Vdd.n570 188.988
R1408 Vdd.n582 Vdd.n576 188.988
R1409 Vdd.n576 Vdd.n569 188.988
R1410 Vdd.n513 Vdd.n494 188.988
R1411 Vdd.n508 Vdd.n494 188.988
R1412 Vdd.n506 Vdd.n500 188.988
R1413 Vdd.n500 Vdd.n493 188.988
R1414 Vdd.n547 Vdd.n539 188.988
R1415 Vdd.n553 Vdd.n547 188.988
R1416 Vdd.n560 Vdd.n541 188.988
R1417 Vdd.n555 Vdd.n541 188.988
R1418 Vdd.n438 Vdd.n419 188.988
R1419 Vdd.n433 Vdd.n419 188.988
R1420 Vdd.n431 Vdd.n425 188.988
R1421 Vdd.n425 Vdd.n418 188.988
R1422 Vdd.n472 Vdd.n464 188.988
R1423 Vdd.n478 Vdd.n472 188.988
R1424 Vdd.n485 Vdd.n466 188.988
R1425 Vdd.n480 Vdd.n466 188.988
R1426 Vdd.n140 Vdd.n139 188.643
R1427 Vdd.n154 Vdd.n153 188.643
R1428 Vdd.n180 Vdd.n179 188.643
R1429 Vdd.n192 Vdd.n191 188.643
R1430 Vdd.n167 Vdd.n166 188.643
R1431 Vdd.n127 Vdd.n126 188.643
R1432 Vdd.n98 Vdd.n97 188.643
R1433 Vdd.n112 Vdd.n111 188.643
R1434 Vdd.n47 Vdd.n35 185.225
R1435 Vdd.n78 Vdd.n35 185.225
R1436 Vdd.n78 Vdd.n77 185.225
R1437 Vdd.n70 Vdd.n69 185.225
R1438 Vdd.n69 Vdd.n49 185.225
R1439 Vdd.n65 Vdd.n49 185.225
R1440 Vdd.n58 Vdd.n57 185.225
R1441 Vdd.n57 Vdd.n52 185.225
R1442 Vdd.n255 Vdd.n254 185.19
R1443 Vdd.n65 Vdd.n64 178.825
R1444 Vdd.n26 Vdd.n25 177.984
R1445 Vdd.n77 Vdd.n36 175.812
R1446 Vdd.n82 Vdd.n81 168.564
R1447 Vdd.n81 Vdd.n32 168.564
R1448 Vdd.n73 Vdd.n32 168.564
R1449 Vdd.n73 Vdd.n41 168.564
R1450 Vdd.n61 Vdd.n41 168.564
R1451 Vdd.n61 Vdd.n54 168.564
R1452 Vdd.n242 Vdd.n205 163.766
R1453 Vdd.n384 Vdd.n348 150.213
R1454 Vdd.n378 Vdd.n377 150.213
R1455 Vdd.n334 Vdd.n333 150.213
R1456 Vdd.n340 Vdd.n304 150.213
R1457 Vdd.n243 Vdd.n201 150.213
R1458 Vdd.n203 Vdd.n201 150.213
R1459 Vdd.n288 Vdd.n287 150.213
R1460 Vdd.n294 Vdd.n258 150.213
R1461 Vdd.n272 Vdd.n271 150.213
R1462 Vdd.n271 Vdd.n259 150.213
R1463 Vdd.n278 Vdd.n259 150.213
R1464 Vdd.n318 Vdd.n317 150.213
R1465 Vdd.n317 Vdd.n305 150.213
R1466 Vdd.n324 Vdd.n305 150.213
R1467 Vdd.n362 Vdd.n361 150.213
R1468 Vdd.n361 Vdd.n349 150.213
R1469 Vdd.n368 Vdd.n349 150.213
R1470 Vdd.n227 Vdd.n226 148.24
R1471 Vdd.n278 Vdd.n169 147.953
R1472 Vdd.n324 Vdd.n143 147.953
R1473 Vdd.n368 Vdd.n116 147.953
R1474 Vdd.n9 Vdd.n1 147.577
R1475 Vdd.n4 Vdd.n1 147.577
R1476 Vdd.n4 Vdd.n0 147.577
R1477 Vdd.n36 Vdd.n27 137.322
R1478 Vdd.n64 Vdd.n63 134.698
R1479 Vdd.n51 Vdd.n39 133.239
R1480 Vdd.n47 Vdd.n46 132.142
R1481 Vdd.n79 Vdd.n26 132.142
R1482 Vdd.n79 Vdd.n78 132.142
R1483 Vdd.n78 Vdd.n34 132.142
R1484 Vdd.n49 Vdd.n34 132.142
R1485 Vdd.n71 Vdd.n47 132.142
R1486 Vdd.n71 Vdd.n70 132.142
R1487 Vdd.n70 Vdd.n48 132.142
R1488 Vdd.n56 Vdd.n49 132.142
R1489 Vdd.n57 Vdd.n56 132.142
R1490 Vdd.n216 Vdd.n215 125.311
R1491 Vdd.n39 Vdd.n38 124.326
R1492 Vdd.n364 Vdd.n100 115.291
R1493 Vdd.n320 Vdd.n129 115.291
R1494 Vdd.n274 Vdd.n156 115.291
R1495 Vdd.n753 Vdd.n740 114.072
R1496 Vdd.n753 Vdd.n752 114.072
R1497 Vdd.n746 Vdd.n745 114.072
R1498 Vdd.n734 Vdd.n733 114.072
R1499 Vdd.n659 Vdd.n658 114.072
R1500 Vdd.n660 Vdd.n659 114.072
R1501 Vdd.n666 Vdd.n645 114.072
R1502 Vdd.n666 Vdd.n665 114.072
R1503 Vdd.n682 Vdd.n681 114.072
R1504 Vdd.n683 Vdd.n682 114.072
R1505 Vdd.n706 Vdd.n705 114.072
R1506 Vdd.n707 Vdd.n706 114.072
R1507 Vdd.n630 Vdd.n629 114.072
R1508 Vdd.n631 Vdd.n630 114.072
R1509 Vdd.n583 Vdd.n582 114.072
R1510 Vdd.n584 Vdd.n583 114.072
R1511 Vdd.n590 Vdd.n569 114.072
R1512 Vdd.n590 Vdd.n589 114.072
R1513 Vdd.n606 Vdd.n605 114.072
R1514 Vdd.n607 Vdd.n606 114.072
R1515 Vdd.n507 Vdd.n506 114.072
R1516 Vdd.n508 Vdd.n507 114.072
R1517 Vdd.n514 Vdd.n493 114.072
R1518 Vdd.n514 Vdd.n513 114.072
R1519 Vdd.n530 Vdd.n529 114.072
R1520 Vdd.n531 Vdd.n530 114.072
R1521 Vdd.n554 Vdd.n553 114.072
R1522 Vdd.n555 Vdd.n554 114.072
R1523 Vdd.n432 Vdd.n431 114.072
R1524 Vdd.n433 Vdd.n432 114.072
R1525 Vdd.n439 Vdd.n418 114.072
R1526 Vdd.n439 Vdd.n438 114.072
R1527 Vdd.n455 Vdd.n454 114.072
R1528 Vdd.n456 Vdd.n455 114.072
R1529 Vdd.n479 Vdd.n478 114.072
R1530 Vdd.n480 Vdd.n479 114.072
R1531 Vdd.n745 Vdd.n723 113.081
R1532 Vdd.n85 Vdd.n84 112.942
R1533 Vdd.n713 Vdd.n712 112.709
R1534 Vdd.n637 Vdd.n636 112.709
R1535 Vdd.n561 Vdd.n560 112.709
R1536 Vdd.n486 Vdd.n485 112.709
R1537 Vdd.n733 Vdd.n720 112.665
R1538 Vdd.n689 Vdd.n688 112.275
R1539 Vdd.n613 Vdd.n612 112.275
R1540 Vdd.n537 Vdd.n536 112.275
R1541 Vdd.n462 Vdd.n461 112.275
R1542 Vdd.n714 Vdd.n691 111.812
R1543 Vdd.n638 Vdd.n615 111.812
R1544 Vdd.n562 Vdd.n539 111.812
R1545 Vdd.n487 Vdd.n464 111.812
R1546 Vdd.n759 Vdd.n722 111.224
R1547 Vdd.n760 Vdd.n721 109.799
R1548 Vdd.n690 Vdd.n667 109.502
R1549 Vdd.n614 Vdd.n591 109.502
R1550 Vdd.n538 Vdd.n515 109.502
R1551 Vdd.n463 Vdd.n440 109.502
R1552 Vdd.n216 Vdd.n206 108.371
R1553 Vdd.n10 Vdd.n9 97.0582
R1554 Vdd.n295 Vdd.n257 93.8044
R1555 Vdd.n341 Vdd.n303 93.8044
R1556 Vdd.n385 Vdd.n347 93.8044
R1557 Vdd.n244 Vdd.n243 87.3417
R1558 Vdd.n243 Vdd.n195 87.3417
R1559 Vdd.n204 Vdd.n203 87.3417
R1560 Vdd.n203 Vdd.n196 87.3417
R1561 Vdd.n272 Vdd.n265 87.3417
R1562 Vdd.n273 Vdd.n272 87.3417
R1563 Vdd.n294 Vdd.n293 87.3417
R1564 Vdd.n293 Vdd.n259 87.3417
R1565 Vdd.n289 Vdd.n259 87.3417
R1566 Vdd.n289 Vdd.n288 87.3417
R1567 Vdd.n318 Vdd.n311 87.3417
R1568 Vdd.n319 Vdd.n318 87.3417
R1569 Vdd.n340 Vdd.n339 87.3417
R1570 Vdd.n339 Vdd.n305 87.3417
R1571 Vdd.n335 Vdd.n305 87.3417
R1572 Vdd.n335 Vdd.n334 87.3417
R1573 Vdd.n362 Vdd.n355 87.3417
R1574 Vdd.n363 Vdd.n362 87.3417
R1575 Vdd.n384 Vdd.n383 87.3417
R1576 Vdd.n383 Vdd.n349 87.3417
R1577 Vdd.n379 Vdd.n349 87.3417
R1578 Vdd.n379 Vdd.n378 87.3417
R1579 Vdd.n372 Vdd.n116 86.2687
R1580 Vdd.n367 Vdd.n116 86.2687
R1581 Vdd.n323 Vdd.n143 86.2687
R1582 Vdd.n328 Vdd.n143 86.2687
R1583 Vdd.n277 Vdd.n169 86.2687
R1584 Vdd.n282 Vdd.n169 86.2687
R1585 Vdd.n227 Vdd.n217 84.7602
R1586 Vdd.n689 Vdd.n668 78.6829
R1587 Vdd.n682 Vdd.n668 78.6829
R1588 Vdd.n613 Vdd.n592 78.6829
R1589 Vdd.n606 Vdd.n592 78.6829
R1590 Vdd.n537 Vdd.n516 78.6829
R1591 Vdd.n530 Vdd.n516 78.6829
R1592 Vdd.n462 Vdd.n441 78.6829
R1593 Vdd.n455 Vdd.n441 78.6829
R1594 Vdd.n734 Vdd.n729 74.9181
R1595 Vdd.n746 Vdd.n741 74.9181
R1596 Vdd.n747 Vdd.n746 74.9181
R1597 Vdd.n735 Vdd.n734 74.9181
R1598 Vdd.n759 Vdd.n758 74.9181
R1599 Vdd.n754 Vdd.n723 74.9181
R1600 Vdd.n754 Vdd.n753 74.9181
R1601 Vdd.n666 Vdd.n644 74.9181
R1602 Vdd.n659 Vdd.n644 74.9181
R1603 Vdd.n713 Vdd.n692 74.9181
R1604 Vdd.n706 Vdd.n692 74.9181
R1605 Vdd.n637 Vdd.n616 74.9181
R1606 Vdd.n630 Vdd.n616 74.9181
R1607 Vdd.n590 Vdd.n568 74.9181
R1608 Vdd.n583 Vdd.n568 74.9181
R1609 Vdd.n514 Vdd.n492 74.9181
R1610 Vdd.n507 Vdd.n492 74.9181
R1611 Vdd.n561 Vdd.n540 74.9181
R1612 Vdd.n554 Vdd.n540 74.9181
R1613 Vdd.n439 Vdd.n417 74.9181
R1614 Vdd.n432 Vdd.n417 74.9181
R1615 Vdd.n486 Vdd.n465 74.9181
R1616 Vdd.n479 Vdd.n465 74.9181
R1617 Vdd.n244 Vdd.n242 73.7887
R1618 Vdd.n758 Vdd.n723 73.4123
R1619 Vdd.n85 Vdd.n26 68.5181
R1620 Vdd.n135 Vdd.n134 61.6672
R1621 Vdd.n139 Vdd.n138 61.6672
R1622 Vdd.n149 Vdd.n148 61.6672
R1623 Vdd.n153 Vdd.n152 61.6672
R1624 Vdd.n175 Vdd.n174 61.6672
R1625 Vdd.n179 Vdd.n178 61.6672
R1626 Vdd.n187 Vdd.n186 61.6672
R1627 Vdd.n191 Vdd.n190 61.6672
R1628 Vdd.n162 Vdd.n161 61.6672
R1629 Vdd.n166 Vdd.n165 61.6672
R1630 Vdd.n122 Vdd.n121 61.6672
R1631 Vdd.n126 Vdd.n125 61.6672
R1632 Vdd.n93 Vdd.n92 61.6672
R1633 Vdd.n97 Vdd.n96 61.6672
R1634 Vdd.n107 Vdd.n106 61.6672
R1635 Vdd.n111 Vdd.n110 61.6672
R1636 Vdd.n2 Vdd.n1 61.6672
R1637 Vdd.n3 Vdd.n0 61.6672
R1638 Vdd.n21 Vdd.n20 61.3942
R1639 Vdd.n295 Vdd.n294 52.0162
R1640 Vdd.n341 Vdd.n340 52.0162
R1641 Vdd.n385 Vdd.n384 52.0162
R1642 Vdd.n255 Vdd.n195 49.2839
R1643 Vdd.n10 Vdd.n0 47.3641
R1644 Vdd.n738 Vdd.n729 46.2505
R1645 Vdd.n738 Vdd.n737 46.2505
R1646 Vdd.n748 Vdd.n747 46.2505
R1647 Vdd.n749 Vdd.n748 46.2505
R1648 Vdd.n750 Vdd.n741 46.2505
R1649 Vdd.n750 Vdd.n749 46.2505
R1650 Vdd.n736 Vdd.n735 46.2505
R1651 Vdd.n737 Vdd.n736 46.2505
R1652 Vdd.n758 Vdd.n757 46.2505
R1653 Vdd.n757 Vdd.n756 46.2505
R1654 Vdd.n755 Vdd.n754 46.2505
R1655 Vdd.n756 Vdd.n755 46.2505
R1656 Vdd.n650 Vdd.n644 46.2505
R1657 Vdd.n650 Vdd.n649 46.2505
R1658 Vdd.n648 Vdd.n646 46.2505
R1659 Vdd.n653 Vdd.n652 46.2505
R1660 Vdd.n676 Vdd.n675 46.2505
R1661 Vdd.n671 Vdd.n669 46.2505
R1662 Vdd.n673 Vdd.n668 46.2505
R1663 Vdd.n673 Vdd.n672 46.2505
R1664 Vdd.n700 Vdd.n699 46.2505
R1665 Vdd.n695 Vdd.n693 46.2505
R1666 Vdd.n697 Vdd.n692 46.2505
R1667 Vdd.n697 Vdd.n696 46.2505
R1668 Vdd.n624 Vdd.n623 46.2505
R1669 Vdd.n619 Vdd.n617 46.2505
R1670 Vdd.n621 Vdd.n616 46.2505
R1671 Vdd.n621 Vdd.n620 46.2505
R1672 Vdd.n574 Vdd.n568 46.2505
R1673 Vdd.n574 Vdd.n573 46.2505
R1674 Vdd.n572 Vdd.n570 46.2505
R1675 Vdd.n577 Vdd.n576 46.2505
R1676 Vdd.n600 Vdd.n599 46.2505
R1677 Vdd.n595 Vdd.n593 46.2505
R1678 Vdd.n597 Vdd.n592 46.2505
R1679 Vdd.n597 Vdd.n596 46.2505
R1680 Vdd.n498 Vdd.n492 46.2505
R1681 Vdd.n498 Vdd.n497 46.2505
R1682 Vdd.n496 Vdd.n494 46.2505
R1683 Vdd.n501 Vdd.n500 46.2505
R1684 Vdd.n524 Vdd.n523 46.2505
R1685 Vdd.n519 Vdd.n517 46.2505
R1686 Vdd.n521 Vdd.n516 46.2505
R1687 Vdd.n521 Vdd.n520 46.2505
R1688 Vdd.n548 Vdd.n547 46.2505
R1689 Vdd.n543 Vdd.n541 46.2505
R1690 Vdd.n545 Vdd.n540 46.2505
R1691 Vdd.n545 Vdd.n544 46.2505
R1692 Vdd.n423 Vdd.n417 46.2505
R1693 Vdd.n423 Vdd.n422 46.2505
R1694 Vdd.n421 Vdd.n419 46.2505
R1695 Vdd.n426 Vdd.n425 46.2505
R1696 Vdd.n449 Vdd.n448 46.2505
R1697 Vdd.n444 Vdd.n442 46.2505
R1698 Vdd.n446 Vdd.n441 46.2505
R1699 Vdd.n446 Vdd.n445 46.2505
R1700 Vdd.n473 Vdd.n472 46.2505
R1701 Vdd.n468 Vdd.n466 46.2505
R1702 Vdd.n470 Vdd.n465 46.2505
R1703 Vdd.n470 Vdd.n469 46.2505
R1704 Vdd.n9 Vdd.n8 46.2505
R1705 Vdd.n5 Vdd.n4 46.2505
R1706 Vdd.n414 Vdd.n413 40.8314
R1707 Vdd.n375 Vdd.n367 37.0005
R1708 Vdd.n375 Vdd.n374 37.0005
R1709 Vdd.n373 Vdd.n372 37.0005
R1710 Vdd.n374 Vdd.n373 37.0005
R1711 Vdd.n331 Vdd.n323 37.0005
R1712 Vdd.n331 Vdd.n330 37.0005
R1713 Vdd.n329 Vdd.n328 37.0005
R1714 Vdd.n330 Vdd.n329 37.0005
R1715 Vdd.n219 Vdd.n217 37.0005
R1716 Vdd.n220 Vdd.n218 37.0005
R1717 Vdd.n208 Vdd.n206 37.0005
R1718 Vdd.n209 Vdd.n207 37.0005
R1719 Vdd.n245 Vdd.n244 37.0005
R1720 Vdd.n197 Vdd.n195 37.0005
R1721 Vdd.n198 Vdd.n197 37.0005
R1722 Vdd.n251 Vdd.n196 37.0005
R1723 Vdd.n204 Vdd.n199 37.0005
R1724 Vdd.n247 Vdd.n199 37.0005
R1725 Vdd.n238 Vdd.n237 37.0005
R1726 Vdd.n234 Vdd.n233 37.0005
R1727 Vdd.n285 Vdd.n277 37.0005
R1728 Vdd.n285 Vdd.n284 37.0005
R1729 Vdd.n283 Vdd.n282 37.0005
R1730 Vdd.n284 Vdd.n283 37.0005
R1731 Vdd.n268 Vdd.n265 37.0005
R1732 Vdd.n268 Vdd.n267 37.0005
R1733 Vdd.n273 Vdd.n264 37.0005
R1734 Vdd.n267 Vdd.n264 37.0005
R1735 Vdd.n293 Vdd.n292 37.0005
R1736 Vdd.n292 Vdd.n291 37.0005
R1737 Vdd.n290 Vdd.n289 37.0005
R1738 Vdd.n291 Vdd.n290 37.0005
R1739 Vdd.n314 Vdd.n311 37.0005
R1740 Vdd.n314 Vdd.n313 37.0005
R1741 Vdd.n319 Vdd.n310 37.0005
R1742 Vdd.n313 Vdd.n310 37.0005
R1743 Vdd.n339 Vdd.n338 37.0005
R1744 Vdd.n338 Vdd.n337 37.0005
R1745 Vdd.n336 Vdd.n335 37.0005
R1746 Vdd.n337 Vdd.n336 37.0005
R1747 Vdd.n358 Vdd.n355 37.0005
R1748 Vdd.n358 Vdd.n357 37.0005
R1749 Vdd.n363 Vdd.n354 37.0005
R1750 Vdd.n357 Vdd.n354 37.0005
R1751 Vdd.n383 Vdd.n382 37.0005
R1752 Vdd.n382 Vdd.n381 37.0005
R1753 Vdd.n380 Vdd.n379 37.0005
R1754 Vdd.n381 Vdd.n380 37.0005
R1755 Vdd.n20 Vdd.n19 37.0005
R1756 Vdd.n16 Vdd.n15 37.0005
R1757 Vdd.n6 Vdd.n5 33.5287
R1758 Vdd.n8 Vdd.n7 33.5287
R1759 Vdd.n252 Vdd.n251 32.732
R1760 Vdd.n246 Vdd.n245 32.732
R1761 Vdd.n407 Vdd.n405 30.8338
R1762 Vdd.n406 Vdd.n404 30.8338
R1763 Vdd.n403 Vdd.n402 28.5005
R1764 Vdd.n288 Vdd.n156 26.8208
R1765 Vdd.n334 Vdd.n129 26.8208
R1766 Vdd.n378 Vdd.n100 26.8208
R1767 Vdd.n752 Vdd.n751 26.4291
R1768 Vdd.n751 Vdd.n727 26.4291
R1769 Vdd.n740 Vdd.n739 26.4291
R1770 Vdd.n739 Vdd.n726 26.4291
R1771 Vdd.n743 Vdd.n722 26.4291
R1772 Vdd.n743 Vdd.n727 26.4291
R1773 Vdd.n745 Vdd.n744 26.4291
R1774 Vdd.n744 Vdd.n727 26.4291
R1775 Vdd.n733 Vdd.n732 26.4291
R1776 Vdd.n732 Vdd.n726 26.4291
R1777 Vdd.n731 Vdd.n721 26.4291
R1778 Vdd.n731 Vdd.n726 26.4291
R1779 Vdd.n661 Vdd.n660 26.4291
R1780 Vdd.n658 Vdd.n657 26.4291
R1781 Vdd.n657 Vdd.n656 26.4291
R1782 Vdd.n654 Vdd.n645 26.4291
R1783 Vdd.n665 Vdd.n664 26.4291
R1784 Vdd.n664 Vdd.n663 26.4291
R1785 Vdd.n677 Vdd.n667 26.4291
R1786 Vdd.n688 Vdd.n687 26.4291
R1787 Vdd.n687 Vdd.n686 26.4291
R1788 Vdd.n684 Vdd.n683 26.4291
R1789 Vdd.n681 Vdd.n680 26.4291
R1790 Vdd.n680 Vdd.n679 26.4291
R1791 Vdd.n701 Vdd.n691 26.4291
R1792 Vdd.n712 Vdd.n711 26.4291
R1793 Vdd.n711 Vdd.n710 26.4291
R1794 Vdd.n708 Vdd.n707 26.4291
R1795 Vdd.n705 Vdd.n704 26.4291
R1796 Vdd.n704 Vdd.n703 26.4291
R1797 Vdd.n625 Vdd.n615 26.4291
R1798 Vdd.n636 Vdd.n635 26.4291
R1799 Vdd.n635 Vdd.n634 26.4291
R1800 Vdd.n632 Vdd.n631 26.4291
R1801 Vdd.n629 Vdd.n628 26.4291
R1802 Vdd.n628 Vdd.n627 26.4291
R1803 Vdd.n585 Vdd.n584 26.4291
R1804 Vdd.n582 Vdd.n581 26.4291
R1805 Vdd.n581 Vdd.n580 26.4291
R1806 Vdd.n578 Vdd.n569 26.4291
R1807 Vdd.n589 Vdd.n588 26.4291
R1808 Vdd.n588 Vdd.n587 26.4291
R1809 Vdd.n601 Vdd.n591 26.4291
R1810 Vdd.n612 Vdd.n611 26.4291
R1811 Vdd.n611 Vdd.n610 26.4291
R1812 Vdd.n608 Vdd.n607 26.4291
R1813 Vdd.n605 Vdd.n604 26.4291
R1814 Vdd.n604 Vdd.n603 26.4291
R1815 Vdd.n509 Vdd.n508 26.4291
R1816 Vdd.n506 Vdd.n505 26.4291
R1817 Vdd.n505 Vdd.n504 26.4291
R1818 Vdd.n502 Vdd.n493 26.4291
R1819 Vdd.n513 Vdd.n512 26.4291
R1820 Vdd.n512 Vdd.n511 26.4291
R1821 Vdd.n525 Vdd.n515 26.4291
R1822 Vdd.n536 Vdd.n535 26.4291
R1823 Vdd.n535 Vdd.n534 26.4291
R1824 Vdd.n532 Vdd.n531 26.4291
R1825 Vdd.n529 Vdd.n528 26.4291
R1826 Vdd.n528 Vdd.n527 26.4291
R1827 Vdd.n549 Vdd.n539 26.4291
R1828 Vdd.n560 Vdd.n559 26.4291
R1829 Vdd.n559 Vdd.n558 26.4291
R1830 Vdd.n556 Vdd.n555 26.4291
R1831 Vdd.n553 Vdd.n552 26.4291
R1832 Vdd.n552 Vdd.n551 26.4291
R1833 Vdd.n434 Vdd.n433 26.4291
R1834 Vdd.n431 Vdd.n430 26.4291
R1835 Vdd.n430 Vdd.n429 26.4291
R1836 Vdd.n427 Vdd.n418 26.4291
R1837 Vdd.n438 Vdd.n437 26.4291
R1838 Vdd.n437 Vdd.n436 26.4291
R1839 Vdd.n450 Vdd.n440 26.4291
R1840 Vdd.n461 Vdd.n460 26.4291
R1841 Vdd.n460 Vdd.n459 26.4291
R1842 Vdd.n457 Vdd.n456 26.4291
R1843 Vdd.n454 Vdd.n453 26.4291
R1844 Vdd.n453 Vdd.n452 26.4291
R1845 Vdd.n474 Vdd.n464 26.4291
R1846 Vdd.n485 Vdd.n484 26.4291
R1847 Vdd.n484 Vdd.n483 26.4291
R1848 Vdd.n481 Vdd.n480 26.4291
R1849 Vdd.n478 Vdd.n477 26.4291
R1850 Vdd.n477 Vdd.n476 26.4291
R1851 Vdd.n7 Vdd.n6 23.2045
R1852 Vdd.n132 Vdd.n131 23.1255
R1853 Vdd.n136 Vdd.n130 23.1255
R1854 Vdd.n146 Vdd.n145 23.1255
R1855 Vdd.n150 Vdd.n144 23.1255
R1856 Vdd.n172 Vdd.n171 23.1255
R1857 Vdd.n176 Vdd.n170 23.1255
R1858 Vdd.n184 Vdd.n183 23.1255
R1859 Vdd.n188 Vdd.n182 23.1255
R1860 Vdd.n159 Vdd.n158 23.1255
R1861 Vdd.n163 Vdd.n157 23.1255
R1862 Vdd.n119 Vdd.n118 23.1255
R1863 Vdd.n123 Vdd.n117 23.1255
R1864 Vdd.n90 Vdd.n89 23.1255
R1865 Vdd.n94 Vdd.n88 23.1255
R1866 Vdd.n104 Vdd.n103 23.1255
R1867 Vdd.n108 Vdd.n102 23.1255
R1868 Vdd.n29 Vdd.n27 20.5561
R1869 Vdd.n81 Vdd.n29 20.5561
R1870 Vdd.n74 Vdd.n39 20.5561
R1871 Vdd.n74 Vdd.n73 20.5561
R1872 Vdd.n46 Vdd.n31 20.5561
R1873 Vdd.n81 Vdd.n31 20.5561
R1874 Vdd.n80 Vdd.n79 20.5561
R1875 Vdd.n81 Vdd.n80 20.5561
R1876 Vdd.n40 Vdd.n34 20.5561
R1877 Vdd.n73 Vdd.n40 20.5561
R1878 Vdd.n72 Vdd.n71 20.5561
R1879 Vdd.n73 Vdd.n72 20.5561
R1880 Vdd.n60 Vdd.n48 20.5561
R1881 Vdd.n61 Vdd.n60 20.5561
R1882 Vdd.n56 Vdd.n50 20.5561
R1883 Vdd.n61 Vdd.n50 20.5561
R1884 Vdd.n63 Vdd.n62 20.5561
R1885 Vdd.n62 Vdd.n61 20.5561
R1886 Vdd.n685 Vdd.n684 19.9367
R1887 Vdd.n678 Vdd.n677 19.9367
R1888 Vdd.n609 Vdd.n608 19.9367
R1889 Vdd.n602 Vdd.n601 19.9367
R1890 Vdd.n533 Vdd.n532 19.9367
R1891 Vdd.n526 Vdd.n525 19.9367
R1892 Vdd.n458 Vdd.n457 19.9367
R1893 Vdd.n451 Vdd.n450 19.9367
R1894 Vdd.n655 Vdd.n654 19.6798
R1895 Vdd.n662 Vdd.n661 19.6798
R1896 Vdd.n709 Vdd.n708 19.6798
R1897 Vdd.n702 Vdd.n701 19.6798
R1898 Vdd.n633 Vdd.n632 19.6798
R1899 Vdd.n626 Vdd.n625 19.6798
R1900 Vdd.n579 Vdd.n578 19.6798
R1901 Vdd.n586 Vdd.n585 19.6798
R1902 Vdd.n503 Vdd.n502 19.6798
R1903 Vdd.n510 Vdd.n509 19.6798
R1904 Vdd.n557 Vdd.n556 19.6798
R1905 Vdd.n550 Vdd.n549 19.6798
R1906 Vdd.n428 Vdd.n427 19.6798
R1907 Vdd.n435 Vdd.n434 19.6798
R1908 Vdd.n482 Vdd.n481 19.6798
R1909 Vdd.n475 Vdd.n474 19.6798
R1910 Vdd.n715 Vdd.n690 19.2662
R1911 Vdd.n640 Vdd.n614 19.2662
R1912 Vdd.n563 Vdd.n538 19.2662
R1913 Vdd.n488 Vdd.n463 19.2662
R1914 Vdd.n371 Vdd.n348 18.5005
R1915 Vdd.n371 Vdd.n353 18.5005
R1916 Vdd.n365 Vdd.n364 18.5005
R1917 Vdd.n365 Vdd.n352 18.5005
R1918 Vdd.n377 Vdd.n376 18.5005
R1919 Vdd.n376 Vdd.n353 18.5005
R1920 Vdd.n321 Vdd.n320 18.5005
R1921 Vdd.n321 Vdd.n308 18.5005
R1922 Vdd.n333 Vdd.n332 18.5005
R1923 Vdd.n332 Vdd.n309 18.5005
R1924 Vdd.n327 Vdd.n304 18.5005
R1925 Vdd.n327 Vdd.n309 18.5005
R1926 Vdd.n222 Vdd.n221 18.5005
R1927 Vdd.n226 Vdd.n225 18.5005
R1928 Vdd.n211 Vdd.n210 18.5005
R1929 Vdd.n215 Vdd.n214 18.5005
R1930 Vdd.n249 Vdd.n201 18.5005
R1931 Vdd.n249 Vdd.n248 18.5005
R1932 Vdd.n254 Vdd.n253 18.5005
R1933 Vdd.n205 Vdd.n202 18.5005
R1934 Vdd.n235 Vdd.n230 18.5005
R1935 Vdd.n231 Vdd.n229 18.5005
R1936 Vdd.n275 Vdd.n274 18.5005
R1937 Vdd.n275 Vdd.n262 18.5005
R1938 Vdd.n287 Vdd.n286 18.5005
R1939 Vdd.n286 Vdd.n263 18.5005
R1940 Vdd.n281 Vdd.n258 18.5005
R1941 Vdd.n281 Vdd.n263 18.5005
R1942 Vdd.n266 Vdd.n257 18.5005
R1943 Vdd.n266 Vdd.n262 18.5005
R1944 Vdd.n271 Vdd.n270 18.5005
R1945 Vdd.n270 Vdd.n262 18.5005
R1946 Vdd.n279 Vdd.n278 18.5005
R1947 Vdd.n279 Vdd.n263 18.5005
R1948 Vdd.n312 Vdd.n303 18.5005
R1949 Vdd.n312 Vdd.n308 18.5005
R1950 Vdd.n317 Vdd.n316 18.5005
R1951 Vdd.n316 Vdd.n308 18.5005
R1952 Vdd.n325 Vdd.n324 18.5005
R1953 Vdd.n325 Vdd.n309 18.5005
R1954 Vdd.n356 Vdd.n347 18.5005
R1955 Vdd.n356 Vdd.n352 18.5005
R1956 Vdd.n361 Vdd.n360 18.5005
R1957 Vdd.n360 Vdd.n352 18.5005
R1958 Vdd.n369 Vdd.n368 18.5005
R1959 Vdd.n369 Vdd.n353 18.5005
R1960 Vdd.n137 Vdd.n136 16.3581
R1961 Vdd.n133 Vdd.n132 16.3581
R1962 Vdd.n151 Vdd.n150 16.3581
R1963 Vdd.n147 Vdd.n146 16.3581
R1964 Vdd.n177 Vdd.n176 16.3581
R1965 Vdd.n173 Vdd.n172 16.3581
R1966 Vdd.n189 Vdd.n188 16.3581
R1967 Vdd.n185 Vdd.n184 16.3581
R1968 Vdd.n164 Vdd.n163 16.3581
R1969 Vdd.n160 Vdd.n159 16.3581
R1970 Vdd.n124 Vdd.n123 16.3581
R1971 Vdd.n120 Vdd.n119 16.3581
R1972 Vdd.n95 Vdd.n94 16.3581
R1973 Vdd.n91 Vdd.n90 16.3581
R1974 Vdd.n109 Vdd.n108 16.3581
R1975 Vdd.n105 Vdd.n104 16.3581
R1976 Vdd.n84 Vdd.n83 15.4172
R1977 Vdd.n83 Vdd.n82 15.4172
R1978 Vdd.n45 Vdd.n30 15.4172
R1979 Vdd.n82 Vdd.n30 15.4172
R1980 Vdd.n42 Vdd.n35 15.4172
R1981 Vdd.n42 Vdd.n32 15.4172
R1982 Vdd.n77 Vdd.n76 15.4172
R1983 Vdd.n76 Vdd.n32 15.4172
R1984 Vdd.n69 Vdd.n68 15.4172
R1985 Vdd.n68 Vdd.n41 15.4172
R1986 Vdd.n66 Vdd.n65 15.4172
R1987 Vdd.n66 Vdd.n41 15.4172
R1988 Vdd.n53 Vdd.n52 15.4172
R1989 Vdd.n54 Vdd.n53 15.4172
R1990 Vdd.n59 Vdd.n58 15.4172
R1991 Vdd.n59 Vdd.n54 15.4172
R1992 Vdd.n17 Vdd.n12 15.4172
R1993 Vdd.n13 Vdd.n11 15.4172
R1994 Vdd.n225 Vdd.n224 13.8458
R1995 Vdd.n223 Vdd.n222 13.8458
R1996 Vdd.n214 Vdd.n213 13.8458
R1997 Vdd.n212 Vdd.n211 13.8458
R1998 Vdd.n236 Vdd.n235 13.8458
R1999 Vdd.n232 Vdd.n231 13.8458
R2000 Vdd.n414 Vdd.n403 13.3491
R2001 Vdd.n137 Vdd.n133 13.1419
R2002 Vdd.n151 Vdd.n147 13.1419
R2003 Vdd.n177 Vdd.n173 13.1419
R2004 Vdd.n189 Vdd.n185 13.1419
R2005 Vdd.n164 Vdd.n160 13.1419
R2006 Vdd.n124 Vdd.n120 13.1419
R2007 Vdd.n95 Vdd.n91 13.1419
R2008 Vdd.n109 Vdd.n105 13.1419
R2009 Vdd.n228 Vdd.n216 12.3889
R2010 Vdd.n302 Vdd.n156 12.157
R2011 Vdd.n390 Vdd.n100 12.0922
R2012 Vdd.n346 Vdd.n129 12.0833
R2013 Vdd.n386 Vdd.n385 12.0162
R2014 Vdd.n342 Vdd.n341 12.0152
R2015 Vdd.n18 Vdd.n17 11.585
R2016 Vdd.n14 Vdd.n13 11.585
R2017 Vdd.n256 Vdd.n255 11.3402
R2018 Vdd.n763 Vdd.n762 11.151
R2019 Vdd.n715 Vdd.n714 10.8138
R2020 Vdd.n563 Vdd.n562 10.8138
R2021 Vdd.n488 Vdd.n487 10.8138
R2022 Vdd.n86 Vdd.n25 10.6765
R2023 Vdd.n296 Vdd.n295 10.623
R2024 Vdd.n51 Vdd.n24 10.2854
R2025 Vdd.n242 Vdd.n241 10.2082
R2026 Vdd.n716 Vdd.n666 9.99521
R2027 Vdd.n641 Vdd.n590 9.99521
R2028 Vdd.n564 Vdd.n514 9.99521
R2029 Vdd.n489 Vdd.n439 9.99521
R2030 Vdd.n761 Vdd.n720 9.91917
R2031 Vdd.n22 Vdd.n21 9.91786
R2032 Vdd.n388 Vdd.n116 9.8005
R2033 Vdd.n344 Vdd.n143 9.8005
R2034 Vdd.n298 Vdd.n169 9.8005
R2035 Vdd Vdd.n180 9.68229
R2036 Vdd.n23 Vdd.n10 9.6755
R2037 Vdd.n86 Vdd.n85 9.66678
R2038 Vdd.n155 Vdd.n154 9.62854
R2039 Vdd.n193 Vdd.n192 9.6275
R2040 Vdd.n128 Vdd.n127 9.62542
R2041 Vdd.n99 Vdd.n98 9.62292
R2042 Vdd.n168 Vdd.n167 9.61667
R2043 Vdd.n228 Vdd.n227 9.59738
R2044 Vdd.n639 Vdd.n638 9.58824
R2045 Vdd.n142 Vdd.n140 9.54371
R2046 Vdd.n114 Vdd.n112 9.54099
R2047 Vdd.n240 Vdd.n239 9.50696
R2048 Vdd.n38 Vdd.n24 9.39898
R2049 Vdd.n761 Vdd.n760 9.3005
R2050 Vdd.n224 Vdd.n223 9.08191
R2051 Vdd.n213 Vdd.n212 9.08191
R2052 Vdd.n236 Vdd.n232 9.08191
R2053 Vdd.n38 Vdd.n36 8.8386
R2054 Vdd.n239 Vdd.n238 8.42627
R2055 Vdd.n140 Vdd.n130 8.26717
R2056 Vdd.n154 Vdd.n144 8.26717
R2057 Vdd.n180 Vdd.n170 8.26717
R2058 Vdd.n192 Vdd.n182 8.26717
R2059 Vdd.n167 Vdd.n157 8.26717
R2060 Vdd.n127 Vdd.n117 8.26717
R2061 Vdd.n98 Vdd.n88 8.26717
R2062 Vdd.n112 Vdd.n102 8.26717
R2063 Vdd.n767 Vdd.n766 7.71333
R2064 Vdd Vdd.n23 7.70011
R2065 Vdd.n18 Vdd.n14 7.52439
R2066 Vdd.n416 Vdd 7.51851
R2067 Vdd.n663 Vdd.n662 6.45728
R2068 Vdd.n656 Vdd.n655 6.45728
R2069 Vdd.n703 Vdd.n702 6.45728
R2070 Vdd.n710 Vdd.n709 6.45728
R2071 Vdd.n627 Vdd.n626 6.45728
R2072 Vdd.n634 Vdd.n633 6.45728
R2073 Vdd.n587 Vdd.n586 6.45728
R2074 Vdd.n580 Vdd.n579 6.45728
R2075 Vdd.n511 Vdd.n510 6.45728
R2076 Vdd.n504 Vdd.n503 6.45728
R2077 Vdd.n551 Vdd.n550 6.45728
R2078 Vdd.n558 Vdd.n557 6.45728
R2079 Vdd.n436 Vdd.n435 6.45728
R2080 Vdd.n429 Vdd.n428 6.45728
R2081 Vdd.n476 Vdd.n475 6.45728
R2082 Vdd.n483 Vdd.n482 6.45728
R2083 Vdd.n679 Vdd.n678 6.20228
R2084 Vdd.n686 Vdd.n685 6.20228
R2085 Vdd.n603 Vdd.n602 6.20228
R2086 Vdd.n610 Vdd.n609 6.20228
R2087 Vdd.n527 Vdd.n526 6.20228
R2088 Vdd.n534 Vdd.n533 6.20228
R2089 Vdd.n452 Vdd.n451 6.20228
R2090 Vdd.n459 Vdd.n458 6.20228
R2091 Vdd.n567 Vdd.n491 5.56249
R2092 Vdd.n719 Vdd.n643 5.48431
R2093 Vdd.n765 Vdd.n567 5.044
R2094 Vdd.n415 Vdd.n414 4.6505
R2095 Vdd.n399 Vdd.n398 4.24736
R2096 Vdd.n409 Vdd.n408 4.02224
R2097 Vdd.n413 Vdd.n412 4.02224
R2098 Vdd.n247 Vdd.n246 3.72621
R2099 Vdd.n252 Vdd.n198 3.72621
R2100 Vdd.n764 Vdd.n719 3.21496
R2101 Vdd.n45 Vdd.n25 3.2005
R2102 Vdd.n766 Vdd 3.12208
R2103 Vdd.n410 Vdd.n409 3.00097
R2104 Vdd.n412 Vdd.n411 3.00097
R2105 Vdd.n400 Vdd.n392 2.90804
R2106 Vdd.n241 Vdd.n240 2.77237
R2107 Vdd.n194 Vdd.n193 2.67413
R2108 Vdd.n416 Vdd.n415 2.52765
R2109 Vdd.n719 Vdd.n718 2.45913
R2110 Vdd.n567 Vdd.n566 2.4555
R2111 Vdd.n411 Vdd.n410 2.04149
R2112 Vdd.n194 Vdd 1.82672
R2113 Vdd.n297 Vdd.n194 1.772
R2114 Vdd.n766 Vdd.n765 1.75219
R2115 Vdd.n690 Vdd.n689 1.74595
R2116 Vdd.n614 Vdd.n613 1.74595
R2117 Vdd.n538 Vdd.n537 1.74595
R2118 Vdd.n463 Vdd.n462 1.74595
R2119 Vdd.n115 Vdd.n101 1.563
R2120 Vdd.n87 Vdd.n24 1.49771
R2121 Vdd.n298 Vdd.n297 1.39712
R2122 Vdd.n386 Vdd.n346 1.33436
R2123 Vdd.n296 Vdd.n256 1.29145
R2124 Vdd.n301 Vdd.n168 1.27405
R2125 Vdd.n256 Vdd 1.2548
R2126 Vdd.n640 Vdd.n639 1.22366
R2127 Vdd.n389 Vdd.n115 1.10834
R2128 Vdd.n241 Vdd.n228 1.10246
R2129 Vdd.n345 Vdd.n142 1.00705
R2130 Vdd.n401 Vdd.n400 0.979016
R2131 Vdd.n297 Vdd.n296 0.959802
R2132 Vdd.n764 Vdd.n763 0.953895
R2133 Vdd.n763 Vdd 0.948843
R2134 Vdd.n87 Vdd.n86 0.903278
R2135 Vdd.n342 Vdd.n302 0.900662
R2136 Vdd.n760 Vdd.n759 0.835283
R2137 Vdd.n639 Vdd 0.814768
R2138 Vdd.n64 Vdd.n51 0.8005
R2139 Vdd.n23 Vdd.n22 0.788852
R2140 Vdd.n344 Vdd.n343 0.772061
R2141 Vdd.n240 Vdd 0.753625
R2142 Vdd.n302 Vdd.n301 0.715329
R2143 Vdd.n765 Vdd.n764 0.663435
R2144 Vdd.n391 Vdd.n390 0.646523
R2145 Vdd Vdd.n416 0.63528
R2146 Vdd.n399 Vdd.n393 0.617037
R2147 Vdd.n714 Vdd.n713 0.610024
R2148 Vdd.n638 Vdd.n637 0.610024
R2149 Vdd.n562 Vdd.n561 0.610024
R2150 Vdd.n487 Vdd.n486 0.610024
R2151 Vdd.n388 Vdd.n387 0.60895
R2152 Vdd.n345 Vdd 0.510601
R2153 Vdd.n767 Vdd.n87 0.482444
R2154 Vdd.n181 Vdd 0.481269
R2155 Vdd.n346 Vdd.n345 0.474526
R2156 Vdd.n387 Vdd.n128 0.445902
R2157 Vdd.n716 Vdd.n715 0.443952
R2158 Vdd.n641 Vdd.n640 0.443952
R2159 Vdd.n564 Vdd.n563 0.443952
R2160 Vdd.n489 Vdd.n488 0.443952
R2161 Vdd.n101 Vdd 0.438
R2162 Vdd.n389 Vdd 0.407318
R2163 Vdd.n391 Vdd.n99 0.402799
R2164 Vdd.n401 Vdd.n391 0.386295
R2165 Vdd.n390 Vdd.n389 0.382318
R2166 Vdd.n343 Vdd.n155 0.378104
R2167 Vdd.n301 Vdd.n300 0.34797
R2168 Vdd.n723 Vdd.n720 0.337342
R2169 Vdd.n22 Vdd 0.315841
R2170 Vdd.n396 Vdd.n392 0.288578
R2171 Vdd.n141 Vdd 0.284591
R2172 Vdd.n400 Vdd.n399 0.257531
R2173 Vdd.n643 Vdd.n641 0.254071
R2174 Vdd.n402 Vdd.n401 0.223227
R2175 Vdd.n566 Vdd.n564 0.214786
R2176 Vdd.n113 Vdd.n101 0.214786
R2177 Vdd.n491 Vdd.n489 0.190381
R2178 Vdd.n300 Vdd 0.18175
R2179 Vdd.n718 Vdd.n717 0.180262
R2180 Vdd.n762 Vdd.n761 0.157444
R2181 Vdd.n300 Vdd.n299 0.13175
R2182 Vdd.n343 Vdd.n342 0.121421
R2183 Vdd.n387 Vdd.n386 0.112202
R2184 Vdd.n395 Vdd.n393 0.104373
R2185 Vdd.n397 Vdd.n395 0.104373
R2186 Vdd.n718 Vdd.n716 0.10169
R2187 Vdd.n717 Vdd 0.09675
R2188 Vdd.n642 Vdd 0.09675
R2189 Vdd.n565 Vdd 0.09675
R2190 Vdd.n490 Vdd 0.09675
R2191 Vdd.n717 Vdd 0.0921667
R2192 Vdd.n642 Vdd 0.0921667
R2193 Vdd.n565 Vdd 0.0921667
R2194 Vdd.n490 Vdd 0.0921667
R2195 Vdd.n491 Vdd.n490 0.0915714
R2196 Vdd.n566 Vdd.n565 0.0671667
R2197 Vdd.n168 Vdd 0.066125
R2198 Vdd.n99 Vdd 0.059875
R2199 Vdd.n128 Vdd 0.057375
R2200 Vdd Vdd.n767 0.05675
R2201 Vdd.n155 Vdd 0.05425
R2202 Vdd.n762 Vdd 0.052375
R2203 Vdd Vdd.n344 0.052375
R2204 Vdd Vdd.n388 0.0476591
R2205 Vdd.n193 Vdd.n181 0.0392583
R2206 Vdd.n142 Vdd.n141 0.0362143
R2207 Vdd.n113 Vdd 0.0348137
R2208 Vdd.n114 Vdd.n113 0.0299118
R2209 Vdd.n643 Vdd.n642 0.027881
R2210 Vdd.n299 Vdd.n298 0.027375
R2211 Vdd.n141 Vdd 0.0266905
R2212 Vdd.n299 Vdd 0.0255
R2213 Vdd.n101 Vdd 0.0183571
R2214 Vdd.n181 Vdd 0.01675
R2215 Vdd.n115 Vdd.n114 0.0152059
R2216 Vdd.n415 Vdd.n402 0.00561364
R2217 Vdd.n398 Vdd.n394 0.00378947
R0 Vss.n496 Vss.n495 1.02685e+06
R1 Vss.n495 Vss.n92 126542
R2 Vss.n126 Vss.n125 55066
R3 Vss.n498 Vss.n497 37820.3
R4 Vss.n127 Vss.n126 36762
R5 Vss.n473 Vss.n212 31750.8
R6 Vss.n365 Vss.n364 29626.4
R7 Vss.n129 Vss.n111 24759.6
R8 Vss.n130 Vss.n109 24489.5
R9 Vss.n111 Vss.n52 23257.1
R10 Vss.n125 Vss.n124 22268
R11 Vss.n368 Vss.n367 20497.5
R12 Vss.n495 Vss.n494 18408.6
R13 Vss.n474 Vss.n211 16430
R14 Vss.n44 Vss.n39 16173.5
R15 Vss.n314 Vss.n252 15290.7
R16 Vss.n310 Vss.n252 15290.7
R17 Vss.n314 Vss.n253 15290.7
R18 Vss.n310 Vss.n253 15290.7
R19 Vss.n307 Vss.n256 15290.7
R20 Vss.n307 Vss.n257 15290.7
R21 Vss.n303 Vss.n256 15290.7
R22 Vss.n303 Vss.n257 15290.7
R23 Vss.n172 Vss.n94 14897.8
R24 Vss.n532 Vss.n531 14877.3
R25 Vss.n531 Vss.n530 14216.9
R26 Vss.n494 Vss.n173 13150
R27 Vss.n130 Vss.n129 12524.6
R28 Vss.n494 Vss.n493 12194.3
R29 Vss.n111 Vss.n110 11666.7
R30 Vss.n212 Vss.n186 11484.6
R31 Vss.n128 Vss.n127 11339.8
R32 Vss.n37 Vss.n31 10110.8
R33 Vss.n256 Vss.n255 9951.21
R34 Vss.n527 Vss.n526 9699.25
R35 Vss.n475 Vss.n210 9610.43
R36 Vss.n518 Vss.n33 8903.4
R37 Vss.n127 Vss.n124 8714.88
R38 Vss.n110 Vss.n109 8607.64
R39 Vss.n339 Vss.n172 7796.45
R40 Vss.n530 Vss.n529 7610.1
R41 Vss.n367 Vss.n366 7300.5
R42 Vss.n526 Vss.n38 7158.07
R43 Vss.n528 Vss.n36 6787.65
R44 Vss.n527 Vss.n37 6615.8
R45 Vss.n366 Vss.n365 6575.56
R46 Vss.n512 Vss.n39 6243.32
R47 Vss.n476 Vss.n209 5323.74
R48 Vss.n163 Vss.n156 5237.88
R49 Vss.n156 Vss.n154 5237.88
R50 Vss.n163 Vss.n157 5237.88
R51 Vss.n157 Vss.n154 5237.88
R52 Vss.n166 Vss.n96 5237.88
R53 Vss.n166 Vss.n97 5237.88
R54 Vss.n170 Vss.n96 5237.88
R55 Vss.n170 Vss.n97 5237.88
R56 Vss.n73 Vss.n32 5209.34
R57 Vss.n86 Vss.n69 5064.06
R58 Vss.n86 Vss.n70 5064.06
R59 Vss.n90 Vss.n69 5064.06
R60 Vss.n90 Vss.n70 5064.06
R61 Vss.n368 Vss.n316 4876
R62 Vss.n74 Vss.n73 4517
R63 Vss.n473 Vss.n213 4470.04
R64 Vss.n367 Vss.n208 4390.72
R65 Vss.n476 Vss.n475 4065.75
R66 Vss.n129 Vss.n128 3754.66
R67 Vss.n213 Vss.n92 3654.25
R68 Vss.n528 Vss.n527 3612.48
R69 Vss.n497 Vss.n94 3558.74
R70 Vss.n528 Vss.n31 3416.07
R71 Vss.n461 Vss.n214 3262.09
R72 Vss.n465 Vss.n461 3262.09
R73 Vss.n471 Vss.n217 3262.09
R74 Vss.n467 Vss.n217 3262.09
R75 Vss.n201 Vss.n196 3262.09
R76 Vss.n205 Vss.n196 3262.09
R77 Vss.n492 Vss.n175 3262.09
R78 Vss.n492 Vss.n176 3262.09
R79 Vss.n364 Vss.n317 3262.09
R80 Vss.n348 Vss.n335 3262.09
R81 Vss.n349 Vss.n348 3262.09
R82 Vss.n364 Vss.n318 3262.09
R83 Vss.n376 Vss.n250 3262.09
R84 Vss.n374 Vss.n250 3262.09
R85 Vss.n382 Vss.n247 3262.09
R86 Vss.n247 Vss.n245 3262.09
R87 Vss.n128 Vss.n123 3242.05
R88 Vss.n513 Vss.n512 3187.75
R89 Vss.n339 Vss.n173 3163.14
R90 Vss.n351 Vss.n350 3153.05
R91 Vss.n531 Vss.n31 3104.73
R92 Vss.n209 Vss.n186 2871.88
R93 Vss.n412 Vss.n391 2856.5
R94 Vss.n420 Vss.n403 2856.5
R95 Vss.n433 Vss.n393 2856.5
R96 Vss.n425 Vss.n406 2856.5
R97 Vss.n285 Vss.n260 2856.5
R98 Vss.n300 Vss.n262 2856.5
R99 Vss.n279 Vss.n269 2856.5
R100 Vss.n295 Vss.n266 2856.5
R101 Vss.n233 Vss.n223 2810.15
R102 Vss.n453 Vss.n233 2810.15
R103 Vss.n459 Vss.n226 2810.15
R104 Vss.n455 Vss.n226 2810.15
R105 Vss.n480 Vss.n187 2810.15
R106 Vss.n190 Vss.n184 2810.15
R107 Vss.n483 Vss.n184 2810.15
R108 Vss.n481 Vss.n480 2810.15
R109 Vss.n352 Vss.n328 2810.15
R110 Vss.n345 Vss.n326 2810.15
R111 Vss.n355 Vss.n326 2810.15
R112 Vss.n353 Vss.n352 2810.15
R113 Vss.n388 Vss.n385 2810.15
R114 Vss.n385 Vss.n243 2810.15
R115 Vss.n440 Vss.n437 2810.15
R116 Vss.n437 Vss.n390 2810.15
R117 Vss.n493 Vss.n174 2780.18
R118 Vss.n39 Vss.n32 2764.69
R119 Vss.n497 Vss.n496 2598.66
R120 Vss.n125 Vss.n38 2531.02
R121 Vss.n509 Vss.n54 2508.85
R122 Vss.n509 Vss.n55 2508.85
R123 Vss.n151 Vss.n54 2508.85
R124 Vss.n151 Vss.n55 2508.85
R125 Vss.n50 Vss.n41 2508.85
R126 Vss.n45 Vss.n41 2508.85
R127 Vss.n50 Vss.n42 2508.85
R128 Vss.n45 Vss.n42 2508.85
R129 Vss.n524 Vss.n514 2508.85
R130 Vss.n519 Vss.n514 2508.85
R131 Vss.n524 Vss.n515 2508.85
R132 Vss.n519 Vss.n515 2508.85
R133 Vss.n104 Vss.n102 2508.85
R134 Vss.n140 Vss.n104 2508.85
R135 Vss.n141 Vss.n102 2508.85
R136 Vss.n141 Vss.n140 2508.85
R137 Vss.n78 Vss.n75 2508.85
R138 Vss.n83 Vss.n75 2508.85
R139 Vss.n83 Vss.n74 2508.85
R140 Vss.n78 Vss.n74 2508.85
R141 Vss.n65 Vss.n63 2508.85
R142 Vss.n499 Vss.n62 2508.85
R143 Vss.n499 Vss.n63 2508.85
R144 Vss.n131 Vss.n107 2508.85
R145 Vss.n136 Vss.n107 2508.85
R146 Vss.n136 Vss.n106 2508.85
R147 Vss.n131 Vss.n106 2508.85
R148 Vss.n116 Vss.n113 2508.85
R149 Vss.n116 Vss.n114 2508.85
R150 Vss.n121 Vss.n114 2508.85
R151 Vss.n121 Vss.n113 2508.85
R152 Vss.n530 Vss.n32 2416.86
R153 Vss.n124 Vss.n123 2355.14
R154 Vss.n498 Vss.n67 2298.37
R155 Vss.n35 Vss.n29 2219.15
R156 Vss.n533 Vss.n29 2219.15
R157 Vss.n35 Vss.n30 2219.15
R158 Vss.n533 Vss.n30 2219.15
R159 Vss.n478 Vss.n477 2169.31
R160 Vss.n529 Vss.n33 2083.94
R161 Vss.n302 Vss.n301 1996.36
R162 Vss.n369 Vss.n315 1855.73
R163 Vss.n474 Vss.n473 1821.36
R164 Vss.n511 Vss.n52 1765.99
R165 Vss.n216 Vss.n214 1755.62
R166 Vss.n471 Vss.n216 1755.62
R167 Vss.n465 Vss.n222 1755.62
R168 Vss.n467 Vss.n222 1755.62
R169 Vss.n225 Vss.n223 1755.62
R170 Vss.n459 Vss.n225 1755.62
R171 Vss.n453 Vss.n231 1755.62
R172 Vss.n455 Vss.n231 1755.62
R173 Vss.n202 Vss.n201 1755.62
R174 Vss.n202 Vss.n175 1755.62
R175 Vss.n205 Vss.n204 1755.62
R176 Vss.n204 Vss.n176 1755.62
R177 Vss.n189 Vss.n187 1755.62
R178 Vss.n190 Vss.n189 1755.62
R179 Vss.n481 Vss.n183 1755.62
R180 Vss.n483 Vss.n183 1755.62
R181 Vss.n341 Vss.n328 1755.62
R182 Vss.n345 Vss.n341 1755.62
R183 Vss.n353 Vss.n325 1755.62
R184 Vss.n355 Vss.n325 1755.62
R185 Vss.n333 Vss.n317 1755.62
R186 Vss.n335 Vss.n333 1755.62
R187 Vss.n331 Vss.n318 1755.62
R188 Vss.n349 Vss.n331 1755.62
R189 Vss.n376 Vss.n246 1755.62
R190 Vss.n382 Vss.n246 1755.62
R191 Vss.n374 Vss.n372 1755.62
R192 Vss.n372 Vss.n245 1755.62
R193 Vss.n388 Vss.n240 1755.62
R194 Vss.n440 Vss.n240 1755.62
R195 Vss.n243 Vss.n241 1755.62
R196 Vss.n390 Vss.n241 1755.62
R197 Vss.n412 Vss.n411 1755.62
R198 Vss.n411 Vss.n403 1755.62
R199 Vss.n405 Vss.n393 1755.62
R200 Vss.n425 Vss.n405 1755.62
R201 Vss.n429 Vss.n394 1755.62
R202 Vss.n429 Vss.n428 1755.62
R203 Vss.n428 Vss.n427 1755.62
R204 Vss.n427 Vss.n400 1755.62
R205 Vss.n261 Vss.n260 1755.62
R206 Vss.n300 Vss.n261 1755.62
R207 Vss.n279 Vss.n271 1755.62
R208 Vss.n271 Vss.n266 1755.62
R209 Vss.n284 Vss.n283 1755.62
R210 Vss.n283 Vss.n273 1755.62
R211 Vss.n273 Vss.n272 1755.62
R212 Vss.n272 Vss.n267 1755.62
R213 Vss.n435 Vss.n208 1613.76
R214 Vss.n92 Vss.n91 1569.53
R215 Vss.n370 Vss.n369 1547.71
R216 Vss.n221 Vss.n216 1506.47
R217 Vss.n222 Vss.n221 1506.47
R218 Vss.n203 Vss.n202 1506.47
R219 Vss.n204 Vss.n203 1506.47
R220 Vss.n333 Vss.n332 1506.47
R221 Vss.n332 Vss.n331 1506.47
R222 Vss.n371 Vss.n246 1506.47
R223 Vss.n372 Vss.n371 1506.47
R224 Vss.n496 Vss.n172 1453.41
R225 Vss.n497 Vss.n93 1448.86
R226 Vss.n369 Vss.n368 1359.1
R227 Vss.n347 Vss.n339 1269.65
R228 Vss.n232 Vss.n211 1260
R229 Vss.n36 Vss.t8 1248.82
R230 Vss.n532 Vss.t8 1248.82
R231 Vss.n477 Vss.n476 1241.33
R232 Vss.n66 Vss.n65 1221.96
R233 Vss.n479 Vss.n206 1173.44
R234 Vss.n334 Vss.n330 1162.98
R235 Vss.n350 Vss.n330 1162.98
R236 Vss.n126 Vss.n37 1159.56
R237 Vss.n365 Vss.n316 1107.17
R238 Vss.n394 Vss.n391 1100.88
R239 Vss.n428 Vss.n398 1100.88
R240 Vss.n411 Vss.n398 1100.88
R241 Vss.n405 Vss.n399 1100.88
R242 Vss.n428 Vss.n399 1100.88
R243 Vss.n433 Vss.n394 1100.88
R244 Vss.n406 Vss.n400 1100.88
R245 Vss.n420 Vss.n400 1100.88
R246 Vss.n275 Vss.n273 1100.88
R247 Vss.n275 Vss.n261 1100.88
R248 Vss.n285 Vss.n284 1100.88
R249 Vss.n293 Vss.n271 1100.88
R250 Vss.n293 Vss.n273 1100.88
R251 Vss.n284 Vss.n269 1100.88
R252 Vss.n295 Vss.n267 1100.88
R253 Vss.n267 Vss.n262 1100.88
R254 Vss.n230 Vss.n225 1054.53
R255 Vss.n231 Vss.n230 1054.53
R256 Vss.n189 Vss.n188 1054.53
R257 Vss.n188 Vss.n183 1054.53
R258 Vss.n341 Vss.n340 1054.53
R259 Vss.n340 Vss.n325 1054.53
R260 Vss.n443 Vss.n240 1054.53
R261 Vss.n443 Vss.n241 1054.53
R262 Vss.n366 Vss.n207 1045.42
R263 Vss.n51 Vss.n40 1013.37
R264 Vss.n44 Vss.n40 1013.37
R265 Vss.n497 Vss.n171 1012.99
R266 Vss.n477 Vss.n208 1009.91
R267 Vss.n313 Vss.n254 993.506
R268 Vss.n311 Vss.n254 993.506
R269 Vss.n313 Vss.n312 993.506
R270 Vss.n312 Vss.n311 993.506
R271 Vss.n306 Vss.n258 993.506
R272 Vss.n306 Vss.n305 993.506
R273 Vss.n304 Vss.n258 993.506
R274 Vss.n305 Vss.n304 993.506
R275 Vss.n347 Vss.n346 978.433
R276 Vss.n529 Vss.n528 969.86
R277 Vss.n77 Vss.n39 941.581
R278 Vss.n512 Vss.n33 883.251
R279 Vss.n351 Vss.n207 839.696
R280 Vss.n212 Vss.n210 781.832
R281 Vss.n512 Vss.n51 724.582
R282 Vss.n482 Vss.n186 700.915
R283 Vss.n316 Vss.n94 696.184
R284 Vss.n113 Vss.n52 670.13
R285 Vss.n482 Vss.n185 667.379
R286 Vss.n545 Vss.n544 598.812
R287 Vss.n75 Vss.n73 597.461
R288 Vss.n543 Vss.n542 594.303
R289 Vss.n138 Vss.n137 575.808
R290 Vss.n526 Vss.n525 560.862
R291 Vss.n475 Vss.n474 559.295
R292 Vss.n200 Vss.n173 557.812
R293 Vss.n315 Vss.n251 556.121
R294 Vss.n309 Vss.n251 556.121
R295 Vss.n153 Vss.n152 539.981
R296 Vss.n302 Vss.n255 498.481
R297 Vss.n123 Vss.n109 497.327
R298 Vss.n213 Vss.n174 496.341
R299 Vss.n454 Vss.n232 486.647
R300 Vss.n200 Vss.n195 432.812
R301 Vss.n206 Vss.n195 432.812
R302 Vss.n436 Vss.n435 396.014
R303 Vss.n257 Vss.n255 390.062
R304 Vss.n518 Vss.n517 381.149
R305 Vss.n517 Vss.n513 363.375
R306 Vss.n478 Vss.n186 362.5
R307 Vss.n165 Vss.n164 360.69
R308 Vss.n155 Vss.n95 360.69
R309 Vss.n162 Vss.n158 340.329
R310 Vss.n159 Vss.n158 340.329
R311 Vss.n160 Vss.n159 340.329
R312 Vss.n167 Vss.n149 340.329
R313 Vss.n168 Vss.n167 340.329
R314 Vss.n169 Vss.n168 340.329
R315 Vss.n87 Vss.n72 329.036
R316 Vss.n88 Vss.n87 329.036
R317 Vss.n89 Vss.n88 329.036
R318 Vss.n210 Vss.n209 322.31
R319 Vss.n85 Vss.n84 308.134
R320 Vss.n308 Vss.n255 283.308
R321 Vss.n479 Vss.n478 275
R322 Vss.n85 Vss.n68 266.399
R323 Vss.n91 Vss.n68 266.399
R324 Vss.n404 Vss.n211 262.546
R325 Vss.n72 Vss.n71 248.095
R326 Vss.n346 Vss.n327 234.871
R327 Vss.n354 Vss.n327 234.871
R328 Vss.n536 Vss.t9 229.403
R329 Vss.n497 Vss.n92 214.635
R330 Vss.n491 Vss.n490 211.953
R331 Vss.n491 Vss.n177 211.953
R332 Vss.n199 Vss.n197 211.953
R333 Vss.n197 Vss.n179 211.953
R334 Vss.n363 Vss.n319 211.953
R335 Vss.n338 Vss.n337 211.953
R336 Vss.n338 Vss.n321 211.953
R337 Vss.n363 Vss.n362 211.953
R338 Vss.n469 Vss.n468 211.953
R339 Vss.n470 Vss.n469 211.953
R340 Vss.n463 Vss.n462 211.953
R341 Vss.n464 Vss.n463 211.953
R342 Vss.n380 Vss.n379 211.953
R343 Vss.n381 Vss.n380 211.953
R344 Vss.n377 Vss.n249 211.953
R345 Vss.n373 Vss.n249 211.953
R346 Vss.n77 Vss.n73 195.47
R347 Vss.n30 Vss.n27 195
R348 Vss.t8 Vss.n30 195
R349 Vss.n29 Vss.n28 195
R350 Vss.t8 Vss.n29 195
R351 Vss.n79 Vss.n78 195
R352 Vss.n78 Vss.n77 195
R353 Vss.n83 Vss.n82 195
R354 Vss.n84 Vss.n83 195
R355 Vss.n65 Vss.n64 195
R356 Vss.n500 Vss.n499 195
R357 Vss.n499 Vss.n498 195
R358 Vss.n132 Vss.n131 195
R359 Vss.n131 Vss.n130 195
R360 Vss.n115 Vss.n113 195
R361 Vss.n142 Vss.n141 195
R362 Vss.n141 Vss.n93 195
R363 Vss.n104 Vss.n103 195
R364 Vss.n138 Vss.n104 195
R365 Vss.n136 Vss.n135 195
R366 Vss.n137 Vss.n136 195
R367 Vss.n119 Vss.n114 195
R368 Vss.n114 Vss.n105 195
R369 Vss.n522 Vss.n515 195
R370 Vss.n517 Vss.n515 195
R371 Vss.n516 Vss.n514 195
R372 Vss.n517 Vss.n514 195
R373 Vss.n48 Vss.n42 195
R374 Vss.n42 Vss.n40 195
R375 Vss.n43 Vss.n41 195
R376 Vss.n41 Vss.n40 195
R377 Vss.n151 Vss.n57 195
R378 Vss.n152 Vss.n151 195
R379 Vss.n509 Vss.n508 195
R380 Vss.n510 Vss.n509 195
R381 Vss.n466 Vss.n460 192.153
R382 Vss.n375 Vss.n370 189.861
R383 Vss.n375 Vss.n244 189.861
R384 Vss.n383 Vss.n244 189.861
R385 Vss.n442 Vss.n389 189.861
R386 Vss.n442 Vss.n441 189.861
R387 Vss.n441 Vss.n436 189.861
R388 Vss.n434 Vss.n392 189.861
R389 Vss.n402 Vss.n392 189.861
R390 Vss.n426 Vss.n402 189.861
R391 Vss.n426 Vss.n404 189.861
R392 Vss.n162 Vss.n161 187.209
R393 Vss.n413 Vss.n396 185.601
R394 Vss.n421 Vss.n419 185.601
R395 Vss.n424 Vss.n423 185.601
R396 Vss.n432 Vss.n395 185.601
R397 Vss.n287 Vss.n286 185.601
R398 Vss.n299 Vss.n298 185.601
R399 Vss.n296 Vss.n265 185.601
R400 Vss.n281 Vss.n280 185.601
R401 Vss.n484 Vss.n182 182.589
R402 Vss.n191 Vss.n182 182.589
R403 Vss.n194 Vss.n180 182.589
R404 Vss.n194 Vss.n193 182.589
R405 Vss.n356 Vss.n324 182.589
R406 Vss.n344 Vss.n324 182.589
R407 Vss.n329 Vss.n322 182.589
R408 Vss.n342 Vss.n329 182.589
R409 Vss.n457 Vss.n456 182.589
R410 Vss.n458 Vss.n457 182.589
R411 Vss.n452 Vss.n235 182.589
R412 Vss.n235 Vss.n234 182.589
R413 Vss.n438 Vss.n238 182.589
R414 Vss.n439 Vss.n438 182.589
R415 Vss.n387 Vss.n386 182.589
R416 Vss.n386 Vss.n237 182.589
R417 Vss.n149 Vss.n148 179.679
R418 Vss.n110 Vss.n38 172.948
R419 Vss.n213 Vss.n185 171.037
R420 Vss.n49 Vss.n43 163.012
R421 Vss.n46 Vss.n43 163.012
R422 Vss.n49 Vss.n48 163.012
R423 Vss.n523 Vss.n516 163.012
R424 Vss.n520 Vss.n516 163.012
R425 Vss.n523 Vss.n522 163.012
R426 Vss.n79 Vss.n76 163.012
R427 Vss.n80 Vss.n79 163.012
R428 Vss.n82 Vss.n76 163.012
R429 Vss.n64 Vss.n60 163.012
R430 Vss.n64 Vss.n61 163.012
R431 Vss.n500 Vss.n61 163.012
R432 Vss.n508 Vss.n507 163.012
R433 Vss.n508 Vss.n56 163.012
R434 Vss.n57 Vss.n56 163.012
R435 Vss.n133 Vss.n132 163.012
R436 Vss.n135 Vss.n108 163.012
R437 Vss.n132 Vss.n108 163.012
R438 Vss.n117 Vss.n115 163.012
R439 Vss.n120 Vss.n115 163.012
R440 Vss.n120 Vss.n119 163.012
R441 Vss.n103 Vss.n101 163.012
R442 Vss.n103 Vss.n100 163.012
R443 Vss.n142 Vss.n101 163.012
R444 Vss.n169 Vss.n148 154.833
R445 Vss.n161 Vss.n160 147.304
R446 Vss.n534 Vss.n533 146.25
R447 Vss.n533 Vss.n532 146.25
R448 Vss.n35 Vss.n34 146.25
R449 Vss.n36 Vss.n35 146.25
R450 Vss.n170 Vss.n169 146.25
R451 Vss.n171 Vss.n170 146.25
R452 Vss.n167 Vss.n166 146.25
R453 Vss.n166 Vss.n165 146.25
R454 Vss.n160 Vss.n157 146.25
R455 Vss.n157 Vss.n95 146.25
R456 Vss.n158 Vss.n156 146.25
R457 Vss.n156 Vss.n153 146.25
R458 Vss.n423 Vss.n406 146.25
R459 Vss.n406 Vss.n404 146.25
R460 Vss.n408 Vss.n399 146.25
R461 Vss.n402 Vss.n399 146.25
R462 Vss.n410 Vss.n398 146.25
R463 Vss.n402 Vss.n398 146.25
R464 Vss.n421 Vss.n420 146.25
R465 Vss.n420 Vss.n404 146.25
R466 Vss.n396 Vss.n391 146.25
R467 Vss.n434 Vss.n391 146.25
R468 Vss.n433 Vss.n432 146.25
R469 Vss.n434 Vss.n433 146.25
R470 Vss.n444 Vss.n443 146.25
R471 Vss.n443 Vss.n442 146.25
R472 Vss.n438 Vss.n437 146.25
R473 Vss.n437 Vss.n436 146.25
R474 Vss.n386 Vss.n385 146.25
R475 Vss.n385 Vss.n384 146.25
R476 Vss.n352 Vss.n329 146.25
R477 Vss.n352 Vss.n351 146.25
R478 Vss.n340 Vss.n323 146.25
R479 Vss.n340 Vss.n327 146.25
R480 Vss.n326 Vss.n324 146.25
R481 Vss.n327 Vss.n326 146.25
R482 Vss.n480 Vss.n194 146.25
R483 Vss.n480 Vss.n479 146.25
R484 Vss.n188 Vss.n181 146.25
R485 Vss.n188 Vss.n185 146.25
R486 Vss.n184 Vss.n182 146.25
R487 Vss.n185 Vss.n184 146.25
R488 Vss.n230 Vss.n229 146.25
R489 Vss.n230 Vss.n224 146.25
R490 Vss.n457 Vss.n226 146.25
R491 Vss.n226 Vss.n224 146.25
R492 Vss.n235 Vss.n233 146.25
R493 Vss.n233 Vss.n224 146.25
R494 Vss.n286 Vss.n285 146.25
R495 Vss.n285 Vss.n259 146.25
R496 Vss.n296 Vss.n295 146.25
R497 Vss.n295 Vss.n294 146.25
R498 Vss.n298 Vss.n262 146.25
R499 Vss.n262 Vss.n259 146.25
R500 Vss.n281 Vss.n269 146.25
R501 Vss.n294 Vss.n269 146.25
R502 Vss.n293 Vss.n292 146.25
R503 Vss.n294 Vss.n293 146.25
R504 Vss.n276 Vss.n275 146.25
R505 Vss.n275 Vss.n259 146.25
R506 Vss.n48 Vss.n47 145.225
R507 Vss.n522 Vss.n521 145.225
R508 Vss.n82 Vss.n81 145.225
R509 Vss.n501 Vss.n500 145.225
R510 Vss.n506 Vss.n57 145.225
R511 Vss.n135 Vss.n134 145.225
R512 Vss.n119 Vss.n118 145.225
R513 Vss.n143 Vss.n142 145.225
R514 Vss.n34 Vss.n28 144.189
R515 Vss.n534 Vss.n28 144.189
R516 Vss.n34 Vss.n27 144.189
R517 Vss.n152 Vss.n150 135.524
R518 Vss.n139 Vss.n138 133.319
R519 Vss.n139 Vss.n93 133.319
R520 Vss.n473 Vss.n472 124.272
R521 Vss.n80 Vss.n75 117.001
R522 Vss.n76 Vss.n74 117.001
R523 Vss.n63 Vss.n60 117.001
R524 Vss.n67 Vss.n63 117.001
R525 Vss.n62 Vss.n61 117.001
R526 Vss.n140 Vss.n100 117.001
R527 Vss.n140 Vss.n139 117.001
R528 Vss.n102 Vss.n101 117.001
R529 Vss.n139 Vss.n102 117.001
R530 Vss.n133 Vss.n107 117.001
R531 Vss.n112 Vss.n107 117.001
R532 Vss.n108 Vss.n106 117.001
R533 Vss.n112 Vss.n106 117.001
R534 Vss.n121 Vss.n120 117.001
R535 Vss.n122 Vss.n121 117.001
R536 Vss.n520 Vss.n519 117.001
R537 Vss.n519 Vss.n518 117.001
R538 Vss.n524 Vss.n523 117.001
R539 Vss.n525 Vss.n524 117.001
R540 Vss.n46 Vss.n45 117.001
R541 Vss.n45 Vss.n44 117.001
R542 Vss.n50 Vss.n49 117.001
R543 Vss.n51 Vss.n50 117.001
R544 Vss.n507 Vss.n55 117.001
R545 Vss.n150 Vss.n55 117.001
R546 Vss.n56 Vss.n54 117.001
R547 Vss.n150 Vss.n54 117.001
R548 Vss.n117 Vss.n116 117.001
R549 Vss.n116 Vss.n53 117.001
R550 Vss.n199 Vss.n198 114.072
R551 Vss.n198 Vss.n177 114.072
R552 Vss.n193 Vss.n192 114.072
R553 Vss.n192 Vss.n191 114.072
R554 Vss.n343 Vss.n342 114.072
R555 Vss.n344 Vss.n343 114.072
R556 Vss.n336 Vss.n319 114.072
R557 Vss.n337 Vss.n336 114.072
R558 Vss.n462 Vss.n218 114.072
R559 Vss.n470 Vss.n218 114.072
R560 Vss.n234 Vss.n227 114.072
R561 Vss.n458 Vss.n227 114.072
R562 Vss.n378 Vss.n377 114.072
R563 Vss.n381 Vss.n378 114.072
R564 Vss.n387 Vss.n239 114.072
R565 Vss.n439 Vss.n239 114.072
R566 Vss.n422 Vss.n401 114.072
R567 Vss.n407 Vss.n395 114.072
R568 Vss.n424 Vss.n407 114.072
R569 Vss.n431 Vss.n430 114.072
R570 Vss.n297 Vss.n264 114.072
R571 Vss.n282 Vss.n277 114.072
R572 Vss.n280 Vss.n274 114.072
R573 Vss.n274 Vss.n265 114.072
R574 Vss.n384 Vss.n242 114.043
R575 Vss.n409 Vss.n401 113.397
R576 Vss.n291 Vss.n264 113.397
R577 Vss.n490 Vss.n489 113.159
R578 Vss.n489 Vss.n179 113.159
R579 Vss.n361 Vss.n321 113.159
R580 Vss.n362 Vss.n361 113.159
R581 Vss.n468 Vss.n219 113.159
R582 Vss.n464 Vss.n219 113.159
R583 Vss.n379 Vss.n236 113.159
R584 Vss.n373 Vss.n236 113.159
R585 Vss.n485 Vss.n484 112.617
R586 Vss.n357 Vss.n356 112.617
R587 Vss.n456 Vss.n228 112.617
R588 Vss.n445 Vss.n238 112.617
R589 Vss.n419 Vss.n418 112.617
R590 Vss.n299 Vss.n263 112.617
R591 Vss.n486 Vss.n180 111.692
R592 Vss.n358 Vss.n322 111.692
R593 Vss.n452 Vss.n451 111.692
R594 Vss.n446 Vss.n237 111.692
R595 Vss.n430 Vss.n397 111.397
R596 Vss.n290 Vss.n277 111.397
R597 Vss.n417 Vss.n413 106.32
R598 Vss.n288 Vss.n287 106.32
R599 Vss.n112 Vss.n105 99.0809
R600 Vss.n535 Vss.n534 98.5969
R601 Vss.n198 Vss.n178 97.8829
R602 Vss.n336 Vss.n320 97.8829
R603 Vss.n220 Vss.n218 97.8829
R604 Vss.n378 Vss.n248 97.8829
R605 Vss.n90 Vss.n89 97.5005
R606 Vss.n91 Vss.n90 97.5005
R607 Vss.n87 Vss.n86 97.5005
R608 Vss.n86 Vss.n85 97.5005
R609 Vss.n364 Vss.n363 97.5005
R610 Vss.n371 Vss.n248 97.5005
R611 Vss.n371 Vss.n244 97.5005
R612 Vss.n380 Vss.n247 97.5005
R613 Vss.n247 Vss.n242 97.5005
R614 Vss.n250 Vss.n249 97.5005
R615 Vss.n370 Vss.n250 97.5005
R616 Vss.n332 Vss.n320 97.5005
R617 Vss.n332 Vss.n330 97.5005
R618 Vss.n348 Vss.n338 97.5005
R619 Vss.n348 Vss.n347 97.5005
R620 Vss.n203 Vss.n178 97.5005
R621 Vss.n203 Vss.n195 97.5005
R622 Vss.n197 Vss.n196 97.5005
R623 Vss.n196 Vss.n195 97.5005
R624 Vss.n492 Vss.n491 97.5005
R625 Vss.n493 Vss.n492 97.5005
R626 Vss.n221 Vss.n220 97.5005
R627 Vss.n221 Vss.n215 97.5005
R628 Vss.n469 Vss.n217 97.5005
R629 Vss.n217 Vss.n215 97.5005
R630 Vss.n463 Vss.n461 97.5005
R631 Vss.n461 Vss.n215 97.5005
R632 Vss.n472 Vss.n215 96.4245
R633 Vss.n466 Vss.n215 96.4245
R634 Vss.n489 Vss.n178 96.377
R635 Vss.n361 Vss.n320 96.377
R636 Vss.n220 Vss.n219 96.377
R637 Vss.n248 Vss.n236 96.377
R638 Vss.n510 Vss.n53 83.8452
R639 Vss.n430 Vss.n429 83.5719
R640 Vss.n429 Vss.n392 83.5719
R641 Vss.n427 Vss.n401 83.5719
R642 Vss.n427 Vss.n426 83.5719
R643 Vss.n419 Vss.n403 83.5719
R644 Vss.n426 Vss.n403 83.5719
R645 Vss.n413 Vss.n412 83.5719
R646 Vss.n412 Vss.n392 83.5719
R647 Vss.n395 Vss.n393 83.5719
R648 Vss.n393 Vss.n392 83.5719
R649 Vss.n425 Vss.n424 83.5719
R650 Vss.n426 Vss.n425 83.5719
R651 Vss.n390 Vss.n238 83.5719
R652 Vss.n441 Vss.n390 83.5719
R653 Vss.n243 Vss.n237 83.5719
R654 Vss.n389 Vss.n243 83.5719
R655 Vss.n388 Vss.n387 83.5719
R656 Vss.n389 Vss.n388 83.5719
R657 Vss.n440 Vss.n439 83.5719
R658 Vss.n441 Vss.n440 83.5719
R659 Vss.n379 Vss.n245 83.5719
R660 Vss.n383 Vss.n245 83.5719
R661 Vss.n374 Vss.n373 83.5719
R662 Vss.n375 Vss.n374 83.5719
R663 Vss.n377 Vss.n376 83.5719
R664 Vss.n376 Vss.n375 83.5719
R665 Vss.n382 Vss.n381 83.5719
R666 Vss.n383 Vss.n382 83.5719
R667 Vss.n349 Vss.n321 83.5719
R668 Vss.n350 Vss.n349 83.5719
R669 Vss.n362 Vss.n318 83.5719
R670 Vss.n350 Vss.n318 83.5719
R671 Vss.n319 Vss.n317 83.5719
R672 Vss.n334 Vss.n317 83.5719
R673 Vss.n337 Vss.n335 83.5719
R674 Vss.n335 Vss.n334 83.5719
R675 Vss.n356 Vss.n355 83.5719
R676 Vss.n355 Vss.n354 83.5719
R677 Vss.n353 Vss.n322 83.5719
R678 Vss.n354 Vss.n353 83.5719
R679 Vss.n342 Vss.n328 83.5719
R680 Vss.n346 Vss.n328 83.5719
R681 Vss.n345 Vss.n344 83.5719
R682 Vss.n346 Vss.n345 83.5719
R683 Vss.n490 Vss.n176 83.5719
R684 Vss.n206 Vss.n176 83.5719
R685 Vss.n205 Vss.n179 83.5719
R686 Vss.n206 Vss.n205 83.5719
R687 Vss.n201 Vss.n199 83.5719
R688 Vss.n201 Vss.n200 83.5719
R689 Vss.n177 Vss.n175 83.5719
R690 Vss.n200 Vss.n175 83.5719
R691 Vss.n484 Vss.n483 83.5719
R692 Vss.n483 Vss.n482 83.5719
R693 Vss.n481 Vss.n180 83.5719
R694 Vss.n482 Vss.n481 83.5719
R695 Vss.n193 Vss.n187 83.5719
R696 Vss.n187 Vss.n174 83.5719
R697 Vss.n191 Vss.n190 83.5719
R698 Vss.n190 Vss.n174 83.5719
R699 Vss.n456 Vss.n455 83.5719
R700 Vss.n455 Vss.n454 83.5719
R701 Vss.n453 Vss.n452 83.5719
R702 Vss.n454 Vss.n453 83.5719
R703 Vss.n234 Vss.n223 83.5719
R704 Vss.n460 Vss.n223 83.5719
R705 Vss.n459 Vss.n458 83.5719
R706 Vss.n460 Vss.n459 83.5719
R707 Vss.n468 Vss.n467 83.5719
R708 Vss.n467 Vss.n466 83.5719
R709 Vss.n465 Vss.n464 83.5719
R710 Vss.n466 Vss.n465 83.5719
R711 Vss.n462 Vss.n214 83.5719
R712 Vss.n472 Vss.n214 83.5719
R713 Vss.n471 Vss.n470 83.5719
R714 Vss.n472 Vss.n471 83.5719
R715 Vss.n287 Vss.n260 83.5719
R716 Vss.n301 Vss.n260 83.5719
R717 Vss.n300 Vss.n299 83.5719
R718 Vss.n301 Vss.n300 83.5719
R719 Vss.n272 Vss.n264 83.5719
R720 Vss.n272 Vss.n270 83.5719
R721 Vss.n283 Vss.n277 83.5719
R722 Vss.n283 Vss.n270 83.5719
R723 Vss.n280 Vss.n279 83.5719
R724 Vss.n279 Vss.n268 83.5719
R725 Vss.n266 Vss.n265 83.5719
R726 Vss.n268 Vss.n266 83.5719
R727 Vss.n89 Vss.n71 80.9417
R728 Vss.n129 Vss.n122 76.7748
R729 Vss.n384 Vss.n383 75.8194
R730 Vss.n389 Vss.n242 75.8194
R731 Vss.n294 Vss.n268 72.0575
R732 Vss.n294 Vss.n270 72.0575
R733 Vss.n270 Vss.n259 72.0575
R734 Vss.n301 Vss.n259 72.0575
R735 Vss.n410 Vss.n409 71.5299
R736 Vss.n423 Vss.n422 71.5299
R737 Vss.n422 Vss.n421 71.5299
R738 Vss.n408 Vss.n407 71.5299
R739 Vss.n432 Vss.n431 71.5299
R740 Vss.n431 Vss.n396 71.5299
R741 Vss.n286 Vss.n282 71.5299
R742 Vss.n298 Vss.n297 71.5299
R743 Vss.n297 Vss.n296 71.5299
R744 Vss.n282 Vss.n281 71.5299
R745 Vss.n292 Vss.n274 71.5299
R746 Vss.n291 Vss.n276 71.5299
R747 Vss.n409 Vss.n408 70.024
R748 Vss.n292 Vss.n291 70.024
R749 Vss.n460 Vss.n224 69.2726
R750 Vss.n454 Vss.n224 69.2726
R751 Vss.n192 Vss.n181 68.5181
R752 Vss.n343 Vss.n323 68.5181
R753 Vss.n229 Vss.n227 68.5181
R754 Vss.n444 Vss.n239 68.5181
R755 Vss.n544 Vss.t7 68.0124
R756 Vss.n544 Vss.t5 68.0124
R757 Vss.n542 Vss.t3 68.0124
R758 Vss.n542 Vss.t1 68.0124
R759 Vss.n418 Vss.n410 67.7652
R760 Vss.n276 Vss.n263 67.7652
R761 Vss.n485 Vss.n181 64.7534
R762 Vss.n357 Vss.n323 64.7534
R763 Vss.n229 Vss.n228 64.7534
R764 Vss.n445 Vss.n444 64.7534
R765 Vss.n309 Vss.n308 63.9569
R766 Vss.n435 Vss.n434 61.4075
R767 Vss.n66 Vss.n62 57.3409
R768 Vss.n67 Vss.n66 56.9871
R769 Vss.n268 Vss.n232 52.9119
R770 Vss.n150 Vss.n53 51.6784
R771 Vss.n512 Vss.n511 51.6474
R772 Vss.n511 Vss.n510 45.8778
R773 Vss.n88 Vss.n70 39.0005
R774 Vss.n70 Vss.n68 39.0005
R775 Vss.n72 Vss.n69 39.0005
R776 Vss.n69 Vss.n68 39.0005
R777 Vss.n535 Vss.n27 38.738
R778 Vss.n122 Vss.n112 34.2377
R779 Vss.n137 Vss.n105 34.2377
R780 Vss.n168 Vss.n97 30.79
R781 Vss.n155 Vss.n97 30.79
R782 Vss.n149 Vss.n96 30.79
R783 Vss.n155 Vss.n96 30.79
R784 Vss.n159 Vss.n154 30.79
R785 Vss.n164 Vss.n154 30.79
R786 Vss.n163 Vss.n162 30.79
R787 Vss.n164 Vss.n163 30.79
R788 Vss.n478 Vss.n207 28.3267
R789 Vss.n537 Vss.t2 28.2503
R790 Vss.n539 Vss.t4 28.2386
R791 Vss.n538 Vss.t6 28.2332
R792 Vss.n541 Vss.t0 28.1447
R793 Vss.n305 Vss.n257 19.5005
R794 Vss.n258 Vss.n256 19.5005
R795 Vss.n312 Vss.n253 19.5005
R796 Vss.n253 Vss.n251 19.5005
R797 Vss.n254 Vss.n252 19.5005
R798 Vss.n252 Vss.n251 19.5005
R799 Vss.n525 Vss.n513 17.7743
R800 Vss.n311 Vss.n310 13.6052
R801 Vss.n310 Vss.n309 13.6052
R802 Vss.n314 Vss.n313 13.6052
R803 Vss.n315 Vss.n314 13.6052
R804 Vss.n307 Vss.n306 13.6052
R805 Vss.n308 Vss.n307 13.6052
R806 Vss.n304 Vss.n303 13.6052
R807 Vss.n303 Vss.n302 13.6052
R808 Vss.n165 Vss.n153 12.6563
R809 Vss.n164 Vss.n155 12.6563
R810 Vss.n171 Vss.n95 12.6563
R811 Vss.n361 Vss.n360 12.4042
R812 Vss.n489 Vss.n488 12.4042
R813 Vss.n447 Vss.n236 12.4042
R814 Vss.n449 Vss.n219 11.4167
R815 Vss.n488 Vss.n486 9.97389
R816 Vss.n360 Vss.n358 9.97389
R817 Vss.n451 Vss.n450 9.97389
R818 Vss.n447 Vss.n446 9.97389
R819 Vss.n47 Vss 9.97133
R820 Vss.n521 Vss 9.97133
R821 Vss.n81 Vss 9.97133
R822 Vss.n502 Vss.n501 9.91696
R823 Vss.n118 Vss.n98 9.91508
R824 Vss.n134 Vss.n99 9.90633
R825 Vss.n144 Vss.n143 9.90383
R826 Vss.n416 Vss.n397 9.89417
R827 Vss.n290 Vss.n289 9.89417
R828 Vss.n71 Vss.n59 9.67897
R829 Vss.n506 Vss.n505 9.49356
R830 Vss.n47 Vss.n46 9.31815
R831 Vss.n521 Vss.n520 9.31815
R832 Vss.n81 Vss.n80 9.31815
R833 Vss.n501 Vss.n60 9.31815
R834 Vss.n507 Vss.n506 9.31815
R835 Vss.n134 Vss.n133 9.31815
R836 Vss.n118 Vss.n117 9.31815
R837 Vss.n143 Vss.n100 9.31815
R838 Vss.n536 Vss.n535 9.3005
R839 Vss.n148 Vss.n147 9.3005
R840 Vss.n161 Vss.n58 9.3005
R841 Vss.n417 Vss.n416 9.3005
R842 Vss.n289 Vss.n288 9.3005
R843 Vss Vss.n415 8.84314
R844 Vss Vss.n545 7.97472
R845 Vss.n1 Vss 6.2505
R846 Vss.n84 Vss.n73 5.77245
R847 Vss.n545 Vss.n543 5.52391
R848 Vss.n547 Vss.n546 5.01259
R849 Vss.n449 Vss.n448 4.55294
R850 Vss Vss.n0 4.48588
R851 Vss.n418 Vss.n417 4.07323
R852 Vss.n288 Vss.n263 4.07323
R853 Vss.n546 Vss 3.3974
R854 Vss.n503 Vss.n59 2.99409
R855 Vss.n504 Vss.n503 2.96087
R856 Vss.n145 Vss.n99 2.91513
R857 Vss.n549 Vss.n2 2.86589
R858 Vss.n548 Vss.n547 2.60559
R859 Vss.n505 Vss.n504 2.39485
R860 Vss.n415 Vss.n0 2.23673
R861 Vss.n548 Vss.n3 2.11622
R862 Vss.n551 Vss.n550 2.01566
R863 Vss.n359 Vss.n3 1.97005
R864 Vss.n409 Vss.n397 1.68471
R865 Vss.n291 Vss.n290 1.68471
R866 Vss.n146 Vss.n98 1.65587
R867 Vss.n354 Vss.n207 1.18076
R868 Vss.n550 Vss.n549 1.08843
R869 Vss.n539 Vss.n538 1.02031
R870 Vss.n450 Vss.n449 0.988
R871 Vss.n503 Vss.n502 0.895311
R872 Vss.n504 Vss.n58 0.883968
R873 Vss.n540 Vss.n537 0.864359
R874 Vss.n448 Vss.n447 0.749298
R875 Vss.n450 Vss.n2 0.747182
R876 Vss.n549 Vss.n548 0.705852
R877 Vss.n360 Vss.n359 0.694856
R878 Vss.n488 Vss.n487 0.683318
R879 Vss.n547 Vss.n26 0.655658
R880 Vss.n487 Vss.n3 0.584667
R881 Vss.n486 Vss.n485 0.582318
R882 Vss.n358 Vss.n357 0.582318
R883 Vss.n451 Vss.n228 0.582318
R884 Vss.n446 Vss.n445 0.582318
R885 Vss.n546 Vss 0.545272
R886 Vss.n145 Vss.n144 0.482872
R887 Vss.n551 Vss.n0 0.388568
R888 Vss.n543 Vss.n541 0.37498
R889 Vss.n147 Vss.n146 0.371535
R890 Vss.n146 Vss.n145 0.365951
R891 Vss Vss.n536 0.341716
R892 Vss.n416 Vss 0.335604
R893 Vss.n147 Vss.n58 0.328726
R894 Vss.n505 Vss 0.328278
R895 Vss.n550 Vss 0.300007
R897 Vss.n289 Vss.n278 0.218362
R898 Vss.n538 Vss.n537 0.191355
R899 Vss.n540 Vss.n539 0.183214
R923 Vss.n278 Vss 0.12175
R924 Vss.n278 Vss 0.119016
R925 Vss.n541 Vss.n540 0.106082
R926 Vss.n414 Vss 0.1055
R927 Vss.n5 Vss.n4 0.0934929
R928 Vss.n7 Vss.n6 0.0934929
R929 Vss.n10 Vss.n9 0.0934929
R930 Vss.n12 Vss.n11 0.0934929
R931 Vss.n18 Vss.n17 0.0934929
R932 Vss.n8 Vss.n7 0.0931571
R933 Vss.n14 Vss.n13 0.0931571
R934 Vss.n15 Vss.n14 0.0931571
R935 Vss.n16 Vss.n15 0.0931571
R936 Vss.n17 Vss.n16 0.0931571
R937 Vss.n20 Vss.n19 0.0931571
R938 Vss.n21 Vss.n20 0.0931571
R939 Vss.n22 Vss.n21 0.0931571
R940 Vss.n23 Vss.n22 0.0931571
R941 Vss.n24 Vss.n23 0.0931571
R942 Vss.n25 Vss.n24 0.0931571
R943 Vss.n6 Vss.n5 0.0928214
R944 Vss.n9 Vss.n8 0.0928214
R945 Vss.n11 Vss.n10 0.0928214
R946 Vss.n13 Vss.n12 0.0928214
R947 Vss.n19 Vss.n18 0.0928214
R948 Vss.n26 Vss.n25 0.0926914
R949 Vss.n487 Vss 0.0689783
R950 Vss.n144 Vss 0.068
R951 Vss.n448 Vss 0.066125
R952 Vss.n99 Vss 0.0655
R953 Vss.n359 Vss 0.0624565
R954 Vss.n1 Vss 0.0617745
R955 Vss.n98 Vss 0.05675
R956 Vss.n502 Vss 0.054875
R957 Vss.n415 Vss 0.053
R958 Vss.n278 Vss 0.0526845
R959 Vss.n59 Vss 0.04175
R960 Vss Vss.n551 0.0352222
R961 Vss.n415 Vss.n414 0.0293208
R962 Vss.n414 Vss 0.0269831
R963 Vss.n2 Vss.n1 0.00172549
R2319 Vin2.n0 Vin2.t1 289.231
R2320 Vin2.n0 Vin2.t0 236.907
R2321 Vin2.n1 Vin2 10.0616
R2322 Vin2 Vin2.n0 1.60764
R2323 Vin2.n1 Vin2 0.688903
R2324 Vin2 Vin2.n1 0.077375
R2325 Vin1.n0 Vin1.t1 289.231
R2326 Vin1.n0 Vin1.t0 236.907
R2327 Vin1.n1 Vin1 7.60808
R2328 Vin1 Vin1.n0 2.79068
R2329 Vin1.n1 Vin1 0.259725
R2330 Vin1 Vin1.n1 0.0705
R2287 Vr.n0 Vr.t1 35.7443
R2288 Vr.n1 Vr.t0 35.2144
R2289 Vr.n1 Vr 7.95204
R2290 Vr.n2 Vr 7.60476
R2291 Vr Vr.n0 2.24341
R2292 Vr.n2 Vr.n1 0.513943
R2293 Vr.n0 Vr 0.063625
R2294 Vr Vr.n2 0.063625
R2313 Iout1.n0 Iout1 11.3901
R2315 Iout1 Iout1.n0 0.059875
R2316 Iout0.n0 Iout0 12.1914
R2318 Iout0 Iout0.n0 0.0605
R2270 Vref4.n2 Vref4.t1 663.212
R2271 Vref4.n0 Vref4.t7 662.317
R2272 Vref4.n2 Vref4.t5 662.317
R2273 Vref4.n0 Vref4.t3 662.312
R2274 Vref4 Vref4.t9 35.7443
R2275 Vref4 Vref4.t8 35.2258
R2276 Vref4.n0 Vref4.t6 28.3652
R2277 Vref4.n0 Vref4.t4 28.2503
R2278 Vref4.n0 Vref4.t0 28.249
R2279 Vref4.n0 Vref4.t2 28.1466
R2280 Vref4 Vref4.n1 10.1787
R2281 Vref4.n3 Vref4.n0 9.84745
R2282 Vref4 Vref4.n3 8.88722
R2283 Vref4.n3 Vref4.n2 8.44664
R2284 Vref4.n1 Vref4 6.72754
R2285 Vref4 Vref4 6.30925
R2286 Vref4.n1 Vref4 5.17691
R2295 Vin3.n0 Vin3.t1 289.231
R2296 Vin3.n0 Vin3.t0 236.907
R2297 Vin3.n1 Vin3 8.34347
R2298 Vin3 Vin3.n0 1.60764
R2299 Vin3.n1 Vin3 0.574277
R2300 Vin3 Vin3.n1 0.059875
R2303 Vin4.n2 Vin4 6.26089
R2304 Vin4.n3 Vin4.n2 2.02998
R2305 Vin4.n2 Vin4.n0 1.98328
R2306 Vin4.n3 Vin4.n1 0.983714
R2307 Vin4 Vin4.n0 0.1955
R2308 Vin4.n0 Vin4 0.0555
R2309 Vin4 Vin4.n3 0.053
R2310 En En.t0 213.084
R2311 En En 12.8455
C4 Vin2 Vss 2.72556f
C5 Vin4 Vss 1.72641f
C6 Vin3 Vss 3.10499f
C7 Vdd.n719 Vss 2.5992f
C8 Vdd.n762 Vss 2.47741f
C9 Vdd.n763 Vss 3.92422f
C10 Vdd.n764 Vss 3.37153f
C11 Vdd.n765 Vss 4.19996f
C12 Vdd.n766 Vss 6.91348f
C0 Vin1 Vin2 3.59613f
C1 Vin3 Vin2 3.72837f
C2 Vin4 Vin3 3.94954f
C3 Vdd Ibias 1.832363f
C13 Vin1 Vss 6.604211f
C18 Iclass1 Vss 3.637646f
C17 Iclass0 Vss 2.451628f
C24 Iout01 Vss 5.717949f
C33 Iout11 Vss 4.43404f
C14 Vin2 Vss 7.014152f
C15 Iout0 Vss 19.595062f
C16 Ibias Vss 31.787489f
C19 Iout1 Vss 12.417305f
C20 En Vss 6.120355f
C21 Vin4 Vss 6.165711f
C22 Vin3 Vss 7.505621f
C35 Vr Vss 16.597572f
C38 Vref4 Vss 21.359648f
C41 Vdd Vss 0.225905p
C42 Vdac0 Vss 15.958673f
C45 Vdac1 Vss 22.824736f
.ends

* expanding   symbol:  /home/eserlis/bump_final_tt.sym # of pins=6
** sym_path: /home/eserlis/bump_final_tt.sym
** sch_path: /home/eserlis/bump_final_tt.sch
.subckt bump_final_tt Vdd Iout Vr Vin Ibias Vss
*.iopin Vss
*.iopin Vin
*.iopin Vr
*.iopin Ibias
*.iopin Iout
*.iopin Vdd
XM3 Ibias Ibias Vss Vss sky130_fd_pr__nfet_01v8 L=1.6 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 Ibias Vss Vss sky130_fd_pr__nfet_01v8 L=1.6 W=0.4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 Vin net1 Vss sky130_fd_pr__nfet_01v8 L=1.6 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net3 Vr net1 Vss sky130_fd_pr__nfet_01v8 L=1.6 W=1.2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net2 net2 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 net4 net2 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM15 Iout net3 net4 Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM16 net5 net3 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM17 Iout net2 net5 Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 net3 net3 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
C3 Ibias Vss 2.492277f
C4 Vdd Vss 11.941113f
C0 net2 Vss 3.09455f
C1 net3 Vss 3.050788f
.ends

* expanding   symbol:  /home/eserlis/ref_gen_tt.sym # of pins=4
** sym_path: /home/eserlis/ref_gen_tt.sym
** sch_path: /home/eserlis/ref_gen_tt.sch
.subckt ref_gen_tt Vdd En Iout Vss
*.iopin Vdd
*.iopin En
*.iopin Iout
*.iopin Vss
XM17 net1 net1 Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Iout net1 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.0 W=1.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 net1 En Vss Vss sky130_fd_pr__nfet_01v8 L=0.5 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

* expanding   symbol:  /home/eserlis/vol_ref_gen_tt.sym # of pins=6
** sym_path: /home/eserlis/vol_ref_gen_tt.sym
** sch_path: /home/eserlis/vol_ref_gen_tt.sch
.subckt vol_ref_gen_tt Vref2 Vdd Vref1 Vss Vref3 Vref4
*.iopin Vdd
*.iopin Vref1
*.iopin Vss
*.iopin Vref2
*.iopin Vref3
*.iopin Vref4
XM17 net1 net1 Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM2 Vref1 Vref1 net1 Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM1 Vref2 Vref2 Vref1 Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 Vref3 Vref3 Vref2 Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM4 Vref4 Vref4 Vref3 Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM5 Vss Vss Vref4 Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
C0 Vref4 Vdd 1.7721f
C1 Vss Vdd 2.960428f
.ends


* expanding   symbol:  /home/eserlis/dac_tt.sym # of pins=8
** sym_path: /home/eserlis/dac_tt.sym
** sch_path: /home/eserlis/dac_tt.sch
.subckt dac_tt Vdd Vss Vin1 Vin2 Vin3 Vin4 Vout1 Vout2
*.iopin Vdd
*.iopin Vss
*.iopin Vin1
*.iopin Vout1
*.iopin Vout2
*.iopin Vin2
*.iopin Vin3
*.iopin Vin4
XM4 Vg Vg Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=10 m=10
R4 Vss Vout1 sky130_fd_pr__res_generic_po W=1 L=1 m=0.01
R1 Vss Vout2 sky130_fd_pr__res_generic_po W=1 L=1 m=0.01
XM31 Vg Vdd Vss Vss sky130_fd_pr__nfet_01v8 L=0.3 W=5 nf=3 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
x1 Vss Vdd net2 Vin4 inv_layout_tt
XM15 net3 Vg net1 Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM18 Vout1 Vg net3 Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x2 Vss Vdd net4 Vin3 inv_layout_tt
x3 Vss Vdd net5 Vin2 inv_layout_tt
x5 Vss Vdd net6 Vin1 inv_layout_tt
x8 net1 Vg Vdd Vin1 net6 Vout1 Vout2 dac_inside_tt
x9 Vdd net7 Vg Vdd Vin4 net2 Vout1 Vout2 dac_inside_tt_v2
x4 net7 net8 Vg Vdd Vin3 net4 Vout1 Vout2 dac_inside_tt_v2
x6 net8 net1 Vg Vdd Vin2 net5 Vout1 Vout2 dac_inside_tt_v2
C0 Vdd Vg 8.131639f
C1 Vout2 Vout1 4.212881f
C2 Vout2 Vdd 2.034039f
C3 Vout1 Vdd 2.236412f
C4 Vg Vss 18.061052f
C5 Vdd Vss 74.997444f
C6 Vout2 Vss 8.7737f
C8 Vin4 Vss 2.224975f
C9 Vout1 Vss 15.433397f
C40 Vg Vss 17.49483f
C12 Vin2 Vss 2.367895f
C15 Vin1 Vss 2.47878f
C18 Vin3 Vss 2.178461f
.ends


* expanding   symbol:  /home/eserlis/ccm_nmos_tt.sym # of pins=3
** sym_path: /home/eserlis/ccm_nmos_tt.sym
** sch_path: /home/eserlis/ccm_nmos_tt.sch
.subckt ccm_nmos_tt Iin Iout Vss
*.iopin Vss
*.iopin Iin
*.iopin Iout
XM3 net1 net1 Vss Vss sky130_fd_pr__nfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net1 Vss Vss sky130_fd_pr__nfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Iin Iin net1 Vss sky130_fd_pr__nfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Iout Iin net2 Vss sky130_fd_pr__nfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
C1 Iin Vss 2.310607f
.ends


* expanding   symbol:  /home/eserlis/wta_pmos_tt.sym # of pins=7
** sym_path: /home/eserlis/wta_pmos_tt.sym
** sch_path: /home/eserlis/wta_pmos_tt.sch
.subckt wta_pmos_tt Vdd Vss Iout1 Iout2 Iin1 Iin2 Ibias
*.iopin Vdd
*.iopin Vss
*.iopin Iout1
*.iopin Iout2
*.iopin Iin1
*.iopin Iin2
*.iopin Ibias
XM11 Iout1 Iin1 Ibias Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Iin1 Ibias Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 Iout2 Iin2 Ibias Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Iin2 Ibias Vdd Vdd sky130_fd_pr__pfet_01v8 L=1.6 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R2 Vss Iout1 sky130_fd_pr__res_generic_po W=10 L=10 m=0.001
R1 Vss Iout2 sky130_fd_pr__res_generic_po W=10 L=10 m=0.001
C0 Iout1 Vdd 5.981853f
C2 Vss Vdd 14.83183f
C3 Iout2 Vdd 6.784562f
.ends


* expanding   symbol:  /home/eserlis/inv_layout_tt.sym # of pins=4
** sym_path: /home/eserlis/inv_layout_tt.sym
** sch_path: /home/eserlis/inv_layout_tt.sch
.subckt inv_layout_tt Vss Vdd Out In
*.iopin Vdd
*.iopin Vss
*.iopin In
*.iopin Out
XM11 Out In Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Out In Vss Vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
C0 Vdd Vss 2.013124f
.ends


* expanding   symbol:  /home/eserlis/dac_inside_tt.sym # of pins=7
** sym_path: /home/eserlis/dac_inside_tt.sym
** sch_path: /home/eserlis/dac_inside_tt.sch
.subckt dac_inside_tt Vupper Vg Vdd Vin Vindot Vout1 Vout2
*.iopin Vg
*.iopin Vin
*.iopin Vdd
*.iopin Vout1
*.iopin Vout2
*.iopin Vupper
*.iopin Vindot
XM8 net1 Vg Vupper Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vout2 Vindot net1 Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout1 Vin net1 Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/eserlis/dac_inside_tt_v2.sym # of pins=8
** sym_path: /home/eserlis/dac_inside_tt_v2.sym
** sch_path: /home/eserlis/dac_inside_tt_v2.sch
.subckt dac_inside_tt_v2 Vupper Vupper_out Vg Vdd Vin Vindot Vout1 Vout2
*.iopin Vg
*.iopin Vin
*.iopin Vdd
*.iopin Vout1
*.iopin Vout2
*.iopin Vupper
*.iopin Vindot
*.iopin Vupper_out
XM8 net1 Vg Vupper Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Vout2 Vindot net1 Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout1 Vin net1 Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 Vupper_out Vg Vupper Vdd sky130_fd_pr__pfet_01v8 L=0.3 W=5 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends