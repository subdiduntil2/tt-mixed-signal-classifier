magic
tech sky130A
magscale 1 2
timestamp 1755119682
<< viali >>
rect 1474 310 4592 454
rect 4636 14 4678 50
rect 1828 -30 1862 4
rect 3136 -960 3190 -926
rect 3014 -2382 3060 -2348
rect 1990 -3332 2028 -3292
rect 1372 -3740 5546 -3688
<< metal1 >>
rect 4634 486 4698 490
rect 1370 482 4698 486
rect 1216 454 4698 482
rect 1216 310 1474 454
rect 4592 310 4698 454
rect 1216 282 4698 310
rect 1370 276 4698 282
rect 1816 4 1868 276
rect 2088 64 2098 124
rect 2198 64 2208 124
rect 1816 -30 1828 4
rect 1862 -30 1868 4
rect 1286 -500 1350 -182
rect 1518 -292 1558 -114
rect 1816 -208 1868 -30
rect 2118 -158 2166 64
rect 1734 -244 1970 -208
rect 1518 -360 1560 -292
rect 2122 -308 2162 -158
rect 1520 -500 1560 -360
rect 1286 -508 1560 -500
rect 2116 -350 2162 -308
rect 2116 -508 2156 -350
rect 1286 -554 2156 -508
rect 1286 -558 2152 -554
rect 1286 -798 1350 -558
rect 1520 -560 2152 -558
rect 2338 -584 2384 -182
rect 2566 -220 2608 276
rect 2850 172 3622 180
rect 2850 124 4386 172
rect 2558 -304 2568 -220
rect 2628 -304 2638 -220
rect 2334 -628 2676 -584
rect 2620 -684 2676 -628
rect 1284 -1546 1352 -798
rect 2624 -1076 2670 -684
rect 2850 -910 2906 124
rect 3606 120 4386 124
rect 3406 -164 3416 -58
rect 3538 -164 3548 -58
rect 4334 -130 4378 120
rect 4594 50 4700 276
rect 4594 14 4636 50
rect 4678 14 4700 50
rect 3092 -336 3102 -226
rect 3236 -336 3246 -226
rect 2852 -992 2900 -910
rect 3114 -926 3224 -336
rect 3114 -960 3136 -926
rect 3190 -960 3224 -926
rect 2626 -1210 2668 -1076
rect 2850 -1298 2902 -992
rect 3114 -1004 3224 -960
rect 3436 -1048 3492 -164
rect 4106 -478 4164 -132
rect 4336 -274 4376 -130
rect 4594 -166 4700 14
rect 4532 -224 4764 -166
rect 4332 -400 4384 -274
rect 4936 -312 4976 -66
rect 4944 -400 4972 -312
rect 4332 -412 4976 -400
rect 5150 -412 5204 -156
rect 4332 -458 5204 -412
rect 4974 -470 5204 -458
rect 4106 -512 4160 -478
rect 3652 -568 4160 -512
rect 3652 -942 3716 -568
rect 5150 -668 5204 -470
rect 5150 -772 5208 -668
rect 3046 -1192 3264 -1156
rect 2848 -1316 2902 -1298
rect 3124 -1478 3178 -1192
rect 3434 -1316 3498 -1048
rect 3654 -1222 3716 -942
rect 5154 -1254 5208 -772
rect 1288 -1614 1352 -1546
rect 1288 -1642 2540 -1614
rect 1288 -1656 2542 -1642
rect 1288 -1658 1352 -1656
rect 2058 -2076 2258 -1876
rect 2506 -2042 2542 -1656
rect 3064 -1678 3264 -1478
rect 5154 -1710 5210 -1254
rect 3530 -1740 5210 -1710
rect 3528 -1766 5210 -1740
rect 2112 -2340 2180 -2076
rect 2712 -2226 2762 -1918
rect 3004 -2040 3064 -2036
rect 2918 -2116 3154 -2040
rect 2712 -2262 2764 -2226
rect 2720 -2340 2764 -2262
rect 2112 -2384 2768 -2340
rect 2122 -2390 2768 -2384
rect 2922 -2584 2954 -2116
rect 3004 -2348 3078 -2326
rect 3004 -2382 3014 -2348
rect 3060 -2382 3078 -2348
rect 3004 -2574 3078 -2382
rect 2860 -2602 2870 -2584
rect 2498 -2654 2870 -2602
rect 2952 -2654 2962 -2584
rect 2498 -2656 2954 -2654
rect 986 -2800 1186 -2704
rect 986 -2804 1338 -2800
rect 1872 -2804 2186 -2802
rect 986 -2806 1576 -2804
rect 1650 -2806 2340 -2804
rect 986 -2856 2340 -2806
rect 986 -2858 1338 -2856
rect 986 -2904 1186 -2858
rect 1478 -2876 2340 -2856
rect 1478 -2880 1800 -2876
rect 1478 -3132 1518 -2880
rect 1656 -3226 1728 -2880
rect 1898 -3130 2122 -3096
rect 1664 -3244 1722 -3226
rect 1982 -3292 2044 -3130
rect 2266 -3146 2338 -2876
rect 2504 -3142 2580 -2656
rect 2266 -3226 2342 -3146
rect 2284 -3244 2342 -3226
rect 1982 -3332 1990 -3292
rect 2028 -3332 2044 -3292
rect 1096 -3646 1296 -3602
rect 1982 -3646 2044 -3332
rect 3002 -3646 3078 -2574
rect 3122 -2602 3154 -2116
rect 3308 -2212 3358 -1930
rect 3528 -2140 3564 -1766
rect 5154 -1770 5210 -1766
rect 3888 -2110 4088 -1910
rect 3308 -2274 3360 -2212
rect 3314 -2394 3360 -2274
rect 3952 -2256 4026 -2110
rect 3952 -2394 4028 -2256
rect 3314 -2452 4028 -2394
rect 3952 -2460 4028 -2452
rect 3106 -2670 3116 -2602
rect 3176 -2670 3186 -2602
rect 1096 -3688 5584 -3646
rect 1096 -3740 1372 -3688
rect 5546 -3740 5584 -3688
rect 1096 -3776 5584 -3740
rect 1096 -3802 1296 -3776
<< via1 >>
rect 2098 64 2198 124
rect 2568 -304 2628 -220
rect 3416 -164 3538 -58
rect 3102 -336 3236 -226
rect 2870 -2654 2952 -2584
rect 3116 -2670 3176 -2602
<< metal2 >>
rect 2098 124 2198 134
rect 2198 80 3496 118
rect 2198 78 3398 80
rect 2098 54 2198 64
rect 3432 -48 3496 80
rect 3416 -58 3538 -48
rect 3416 -174 3538 -164
rect 2568 -220 2628 -210
rect 3102 -226 3236 -216
rect 2628 -300 3102 -228
rect 2568 -314 2628 -304
rect 3102 -346 3236 -336
rect 2870 -2584 2952 -2574
rect 3116 -2602 3176 -2592
rect 2952 -2654 3116 -2608
rect 2870 -2664 2952 -2654
rect 3116 -2680 3176 -2670
use sky130_fd_pr__nfet_01v8_484FDA  XM3
timestamp 1754378775
transform 1 0 1704 0 1 -3120
box -356 -252 356 252
use sky130_fd_pr__nfet_01v8_484FDA  XM4
timestamp 1754378775
transform 1 0 2310 0 1 -3120
box -356 -252 356 252
use sky130_fd_pr__nfet_01v8_7QMDBN  XM5
timestamp 1754378775
transform 1 0 2734 0 1 -2092
box -356 -330 356 330
use sky130_fd_pr__nfet_01v8_7QMDBN  XM6
timestamp 1754378775
transform 1 0 3340 0 1 -2092
box -356 -330 356 330
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM13
timestamp 1754378775
transform 1 0 1542 0 1 -231
box -356 -269 356 269
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM14
timestamp 1754378775
transform 1 0 2148 0 1 -231
box -356 -269 356 269
use sky130_fd_pr__pfet_01v8_Q6Z9BJ  XM15
timestamp 1754378775
transform 1 0 2854 0 1 -1179
box -356 -279 356 279
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM16
timestamp 1754378775
transform 1 0 4352 0 1 -191
box -356 -269 356 269
use sky130_fd_pr__pfet_01v8_Q6Z9BJ  XM17
timestamp 1754378775
transform 1 0 3460 0 1 -1179
box -356 -279 356 279
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM18
timestamp 1754378775
transform 1 0 4958 0 1 -191
box -356 -269 356 269
<< labels >>
flabel metal1 2058 -2076 2258 -1876 0 FreeSans 256 0 0 0 Vin
port 3 nsew
flabel metal1 3888 -2110 4088 -1910 0 FreeSans 256 0 0 0 Vr
port 2 nsew
flabel metal1 1096 -3802 1296 -3602 0 FreeSans 256 0 0 0 Vss
port 5 nsew
flabel metal1 1216 282 1416 482 0 FreeSans 256 0 0 0 Vdd
port 0 nsew
flabel metal1 3064 -1678 3264 -1478 0 FreeSans 256 0 0 0 Iout
port 1 nsew
rlabel metal1 1528 -542 1578 -518 1 l3
rlabel metal1 4908 -1758 4958 -1734 1 l4
rlabel metal1 2430 -616 2480 -592 1 l5
rlabel metal1 3752 -556 3802 -532 1 l6
flabel metal1 986 -2904 1186 -2704 0 FreeSans 256 0 0 0 Ibias
port 4 nsew
<< end >>
