magic
tech sky130A
magscale 1 2
timestamp 1755355673
<< locali >>
rect 152 580 2628 614
rect 152 514 280 580
rect 2606 514 2628 580
rect 152 506 2628 514
rect 392 -2186 2776 -2164
rect 392 -2258 544 -2186
rect 2742 -2258 2776 -2186
rect 392 -2268 2776 -2258
<< viali >>
rect 280 514 2606 580
rect 1448 236 1492 272
rect 2118 246 2154 280
rect 662 -566 698 -474
rect 642 -1262 686 -1186
rect 544 -2258 2742 -2186
<< metal1 >>
rect 22 614 222 656
rect 22 590 2628 614
rect 22 580 2630 590
rect 22 514 280 580
rect 2606 530 2630 580
rect 2606 514 2628 530
rect 22 506 2628 514
rect 22 456 222 506
rect 542 380 616 506
rect 1114 458 1226 506
rect 536 -442 616 380
rect 1102 370 1112 458
rect 1234 370 1244 458
rect 1428 308 1514 506
rect 1422 296 1514 308
rect 1422 272 1520 296
rect 1422 246 1448 272
rect 1424 236 1448 246
rect 1492 236 1520 272
rect 1424 234 1520 236
rect 2110 280 2160 506
rect 2110 246 2118 280
rect 2154 246 2160 280
rect 1424 230 1516 234
rect 2110 230 2160 246
rect 718 -6 784 82
rect 716 -50 784 -6
rect 716 -194 780 -50
rect 934 -82 984 140
rect 1128 0 1138 76
rect 1194 0 1204 76
rect 1318 -50 1368 142
rect 1920 60 1980 156
rect 2112 60 2122 90
rect 940 -86 978 -82
rect 938 -156 978 -86
rect 1066 -88 1374 -50
rect 1542 -56 1584 58
rect 1404 -88 1584 -56
rect 1326 -156 1364 -88
rect 940 -166 978 -156
rect 922 -178 978 -166
rect 716 -250 782 -194
rect 716 -316 748 -250
rect 738 -322 748 -316
rect 818 -322 828 -250
rect 922 -388 972 -178
rect 1088 -194 1396 -156
rect 1132 -314 1142 -234
rect 1196 -314 1206 -234
rect 1080 -404 1120 -376
rect 1212 -384 1268 -376
rect 1212 -404 1290 -384
rect 1326 -392 1376 -194
rect 1542 -232 1584 -88
rect 1490 -330 1500 -232
rect 1584 -330 1594 -232
rect 1706 -236 1774 52
rect 1920 26 2122 60
rect 1920 8 1980 26
rect 1916 -80 1980 8
rect 2112 2 2122 26
rect 2186 2 2196 90
rect 1916 -168 1962 -80
rect 2100 -88 2240 -48
rect 2302 -72 2362 164
rect 1706 -304 1744 -236
rect 1734 -324 1744 -304
rect 1808 -324 1818 -236
rect 1906 -404 1966 -168
rect 2108 -198 2248 -158
rect 2316 -168 2362 -72
rect 2108 -328 2118 -240
rect 2182 -328 2192 -240
rect 2306 -404 2366 -168
rect 2532 -238 2600 52
rect 2490 -324 2500 -238
rect 2564 -304 2600 -238
rect 2564 -324 2574 -304
rect 536 -474 724 -442
rect 2758 -450 2958 -390
rect 2138 -456 2958 -450
rect 536 -566 662 -474
rect 698 -566 724 -474
rect 2114 -526 2124 -456
rect 2176 -526 2958 -456
rect 2138 -532 2958 -526
rect 536 -574 724 -566
rect 536 -610 610 -574
rect 686 -576 724 -574
rect 532 -664 612 -610
rect 530 -1162 614 -664
rect 732 -982 784 -674
rect 940 -826 986 -590
rect 1328 -606 1374 -572
rect 2758 -590 2958 -532
rect 1132 -734 1142 -658
rect 1194 -734 1204 -658
rect 1314 -674 1374 -606
rect 1938 -592 1958 -590
rect 1542 -674 1594 -666
rect 1938 -670 1986 -592
rect 2110 -670 2120 -666
rect 1314 -724 1594 -674
rect 1314 -786 1374 -724
rect 1012 -820 1394 -786
rect 946 -900 980 -826
rect 1326 -892 1360 -820
rect 732 -1052 760 -982
rect 814 -1052 824 -982
rect 732 -1054 784 -1052
rect 942 -1136 988 -900
rect 1026 -926 1408 -892
rect 1134 -1054 1144 -978
rect 1196 -1054 1206 -978
rect 1322 -1136 1368 -926
rect 1542 -982 1594 -724
rect 1744 -980 1772 -674
rect 1938 -706 2120 -670
rect 1934 -722 2120 -706
rect 1934 -916 1988 -722
rect 2110 -744 2120 -722
rect 2174 -744 2184 -666
rect 2308 -784 2350 -602
rect 2012 -816 2364 -784
rect 1932 -928 1988 -916
rect 1506 -1052 1516 -982
rect 1570 -1046 1594 -982
rect 1570 -1052 1580 -1046
rect 1740 -1050 1750 -980
rect 1804 -1050 1814 -980
rect 1932 -1110 1974 -928
rect 2080 -932 2266 -892
rect 2316 -926 2350 -816
rect 2114 -1060 2124 -982
rect 2178 -1060 2188 -982
rect 1932 -1114 2296 -1110
rect 1944 -1142 2296 -1114
rect 2314 -1124 2356 -926
rect 2528 -984 2556 -692
rect 2494 -1054 2504 -984
rect 2558 -992 2568 -984
rect 2754 -992 2952 -918
rect 2558 -1038 2952 -992
rect 2558 -1054 2568 -1038
rect 2754 -1118 2952 -1038
rect 526 -1186 724 -1162
rect 526 -1262 642 -1186
rect 686 -1262 724 -1186
rect 2098 -1254 2108 -1194
rect 2172 -1204 2182 -1194
rect 2768 -1204 2968 -1176
rect 2172 -1250 2968 -1204
rect 2172 -1254 2182 -1250
rect 526 -1282 724 -1262
rect 742 -1708 780 -1414
rect 936 -1454 1000 -1318
rect 936 -1550 1002 -1454
rect 1124 -1484 1134 -1382
rect 1194 -1484 1204 -1382
rect 1312 -1408 1376 -1306
rect 1312 -1462 1538 -1408
rect 942 -1620 1002 -1550
rect 1094 -1560 1280 -1520
rect 1312 -1538 1376 -1462
rect 742 -1796 752 -1708
rect 820 -1796 830 -1708
rect 940 -1852 1004 -1620
rect 1084 -1668 1270 -1628
rect 1314 -1634 1374 -1538
rect 1314 -1680 1382 -1634
rect 1126 -1804 1136 -1702
rect 1196 -1804 1206 -1702
rect 1318 -1866 1382 -1680
rect 1542 -1712 1580 -1404
rect 1934 -1406 1998 -1318
rect 2114 -1406 2124 -1396
rect 1732 -1702 1770 -1418
rect 1934 -1460 2124 -1406
rect 1934 -1550 1998 -1460
rect 2114 -1468 2124 -1460
rect 2182 -1468 2192 -1396
rect 1936 -1632 1996 -1550
rect 2086 -1560 2272 -1520
rect 2306 -1564 2370 -1332
rect 2768 -1376 2968 -1250
rect 1936 -1672 2004 -1632
rect 2090 -1672 2276 -1632
rect 2310 -1644 2370 -1564
rect 1506 -1792 1516 -1712
rect 1580 -1792 1590 -1712
rect 1732 -1794 1748 -1702
rect 1806 -1794 1816 -1702
rect 1940 -1864 2004 -1672
rect 2108 -1784 2118 -1712
rect 2176 -1784 2186 -1712
rect 2298 -1878 2362 -1646
rect 2534 -1702 2572 -1408
rect 2494 -1794 2504 -1702
rect 2562 -1722 2572 -1702
rect 2740 -1722 2940 -1648
rect 2562 -1790 2940 -1722
rect 2562 -1794 2572 -1790
rect 2740 -1848 2940 -1790
rect 2098 -2114 2108 -2044
rect 2200 -2114 2210 -2044
rect 316 -2126 394 -2118
rect 262 -2164 462 -2126
rect 2120 -2164 2168 -2114
rect 262 -2186 2776 -2164
rect 262 -2258 544 -2186
rect 2742 -2258 2776 -2186
rect 262 -2268 2776 -2258
rect 262 -2326 462 -2268
<< via1 >>
rect 1112 370 1234 458
rect 1138 0 1194 76
rect 748 -322 818 -250
rect 1142 -314 1196 -234
rect 1500 -330 1584 -232
rect 2122 2 2186 90
rect 1744 -324 1808 -236
rect 2118 -328 2182 -240
rect 2500 -324 2564 -238
rect 2124 -526 2176 -456
rect 1142 -734 1194 -658
rect 760 -1052 814 -982
rect 1144 -1054 1196 -978
rect 2120 -744 2174 -666
rect 1516 -1052 1570 -982
rect 1750 -1050 1804 -980
rect 2124 -1060 2178 -982
rect 2504 -1054 2558 -984
rect 2108 -1254 2172 -1194
rect 1134 -1484 1194 -1382
rect 752 -1796 820 -1708
rect 1136 -1804 1196 -1702
rect 2124 -1468 2182 -1396
rect 1516 -1792 1580 -1712
rect 1748 -1794 1806 -1702
rect 2118 -1784 2176 -1712
rect 2504 -1794 2562 -1702
rect 2108 -2114 2200 -2044
<< metal2 >>
rect 1112 458 1234 468
rect 1112 360 1234 370
rect 1150 86 1212 360
rect 1138 76 1212 86
rect 2122 90 2186 100
rect 1194 30 1212 76
rect 1138 -10 1194 0
rect 2118 2 2122 84
rect 2118 -8 2186 2
rect 744 -230 860 -220
rect 1152 -224 1180 -10
rect 1142 -234 1196 -224
rect 1142 -324 1196 -314
rect 1500 -232 1584 -222
rect 1500 -340 1584 -330
rect 1706 -226 1828 -216
rect 744 -350 860 -340
rect 2118 -230 2178 -8
rect 2470 -216 2592 -206
rect 2118 -240 2182 -230
rect 2118 -338 2182 -328
rect 1706 -362 1828 -352
rect 2128 -446 2160 -338
rect 2470 -352 2592 -342
rect 2124 -456 2176 -446
rect 1146 -526 2124 -456
rect 1146 -528 2176 -526
rect 1146 -570 1186 -528
rect 2124 -536 2176 -528
rect 1148 -648 1178 -570
rect 1142 -658 1194 -648
rect 1142 -744 1194 -734
rect 2120 -666 2174 -656
rect 742 -974 840 -964
rect 1158 -968 1190 -744
rect 2120 -754 2174 -744
rect 1730 -960 1828 -950
rect 1144 -978 1196 -968
rect 1144 -1064 1196 -1054
rect 1502 -972 1600 -962
rect 742 -1082 840 -1072
rect 2134 -972 2162 -754
rect 2482 -968 2580 -958
rect 1730 -1068 1828 -1058
rect 2124 -982 2178 -972
rect 2124 -1070 2178 -1060
rect 1502 -1080 1600 -1070
rect 2130 -1184 2168 -1070
rect 2482 -1076 2580 -1066
rect 2108 -1192 2172 -1184
rect 1140 -1194 2172 -1192
rect 1140 -1250 2108 -1194
rect 1140 -1276 1186 -1250
rect 2108 -1264 2172 -1254
rect 1146 -1372 1186 -1276
rect 1134 -1382 1194 -1372
rect 2124 -1396 2182 -1386
rect 2124 -1478 2182 -1468
rect 1134 -1494 1194 -1484
rect 736 -1696 838 -1686
rect 1144 -1692 1182 -1494
rect 736 -1818 838 -1808
rect 1136 -1702 1196 -1692
rect 1136 -1814 1196 -1804
rect 1502 -1696 1604 -1686
rect 1502 -1818 1604 -1808
rect 1724 -1690 1822 -1680
rect 2134 -1702 2168 -1478
rect 2484 -1684 2582 -1674
rect 2118 -1712 2176 -1702
rect 2118 -1794 2176 -1784
rect 1724 -1820 1822 -1810
rect 2134 -1798 2168 -1794
rect 2134 -2034 2164 -1798
rect 2484 -1814 2582 -1804
rect 2108 -2044 2200 -2034
rect 2108 -2124 2200 -2114
<< via2 >>
rect 744 -250 860 -230
rect 744 -322 748 -250
rect 748 -322 818 -250
rect 818 -322 860 -250
rect 744 -340 860 -322
rect 1500 -330 1584 -232
rect 1706 -236 1828 -226
rect 1706 -324 1744 -236
rect 1744 -324 1808 -236
rect 1808 -324 1828 -236
rect 1706 -352 1828 -324
rect 2470 -238 2592 -216
rect 2470 -324 2500 -238
rect 2500 -324 2564 -238
rect 2564 -324 2592 -238
rect 2470 -342 2592 -324
rect 742 -982 840 -974
rect 742 -1052 760 -982
rect 760 -1052 814 -982
rect 814 -1052 840 -982
rect 742 -1072 840 -1052
rect 1502 -982 1600 -972
rect 1502 -1052 1516 -982
rect 1516 -1052 1570 -982
rect 1570 -1052 1600 -982
rect 1502 -1070 1600 -1052
rect 1730 -980 1828 -960
rect 1730 -1050 1750 -980
rect 1750 -1050 1804 -980
rect 1804 -1050 1828 -980
rect 1730 -1058 1828 -1050
rect 2482 -984 2580 -968
rect 2482 -1054 2504 -984
rect 2504 -1054 2558 -984
rect 2558 -1054 2580 -984
rect 2482 -1066 2580 -1054
rect 736 -1708 838 -1696
rect 736 -1796 752 -1708
rect 752 -1796 820 -1708
rect 820 -1796 838 -1708
rect 736 -1808 838 -1796
rect 1502 -1712 1604 -1696
rect 1502 -1792 1516 -1712
rect 1516 -1792 1580 -1712
rect 1580 -1792 1604 -1712
rect 1502 -1808 1604 -1792
rect 1724 -1702 1822 -1690
rect 2484 -1702 2582 -1684
rect 1724 -1794 1748 -1702
rect 1748 -1794 1806 -1702
rect 1806 -1794 1822 -1702
rect 2484 -1794 2504 -1702
rect 2504 -1794 2562 -1702
rect 2562 -1794 2582 -1702
rect 1724 -1810 1822 -1794
rect 2484 -1804 2582 -1794
<< metal3 >>
rect 2460 -216 2602 -211
rect 734 -230 870 -225
rect 1696 -226 1838 -221
rect 734 -340 744 -230
rect 860 -236 870 -230
rect 1490 -232 1594 -227
rect 1490 -236 1500 -232
rect 860 -296 1500 -236
rect 860 -340 870 -296
rect 1478 -310 1500 -296
rect 1490 -330 1500 -310
rect 1584 -246 1594 -232
rect 1696 -246 1706 -226
rect 1584 -310 1706 -246
rect 1584 -330 1594 -310
rect 1490 -335 1594 -330
rect 734 -345 870 -340
rect 1696 -352 1706 -310
rect 1828 -246 1838 -226
rect 2460 -246 2470 -216
rect 1828 -310 2470 -246
rect 1828 -352 1838 -310
rect 2460 -342 2470 -310
rect 2592 -342 2602 -216
rect 2460 -347 2602 -342
rect 1696 -357 1838 -352
rect 1720 -960 1838 -955
rect 732 -974 850 -969
rect 732 -1072 742 -974
rect 840 -1002 850 -974
rect 1492 -972 1610 -967
rect 1492 -1002 1502 -972
rect 840 -1062 1502 -1002
rect 840 -1072 850 -1062
rect 732 -1077 850 -1072
rect 1492 -1070 1502 -1062
rect 1600 -1002 1610 -972
rect 1720 -1002 1730 -960
rect 1600 -1058 1730 -1002
rect 1828 -1002 1838 -960
rect 2472 -968 2590 -963
rect 2472 -1002 2482 -968
rect 1828 -1058 2482 -1002
rect 1600 -1062 2482 -1058
rect 1600 -1070 1610 -1062
rect 1720 -1063 1838 -1062
rect 1492 -1075 1610 -1070
rect 2472 -1066 2482 -1062
rect 2580 -1066 2590 -968
rect 2472 -1071 2590 -1066
rect 2474 -1684 2592 -1679
rect 1714 -1690 1832 -1685
rect 726 -1696 848 -1691
rect 726 -1808 736 -1696
rect 838 -1720 848 -1696
rect 1492 -1696 1614 -1691
rect 1492 -1720 1502 -1696
rect 838 -1782 1502 -1720
rect 838 -1808 848 -1782
rect 726 -1813 848 -1808
rect 1492 -1808 1502 -1782
rect 1604 -1720 1614 -1696
rect 1714 -1720 1724 -1690
rect 1604 -1782 1724 -1720
rect 1604 -1808 1614 -1782
rect 1492 -1813 1614 -1808
rect 1714 -1810 1724 -1782
rect 1822 -1720 1832 -1690
rect 2474 -1720 2484 -1684
rect 1822 -1782 2484 -1720
rect 1822 -1810 1832 -1782
rect 2474 -1804 2484 -1782
rect 2582 -1804 2592 -1684
rect 2474 -1809 2592 -1804
rect 1714 -1815 1832 -1810
use sky130_fd_pr__pfet_01v8_8WDS2C  XM1
timestamp 1754378775
transform 1 0 1165 0 1 -859
box -545 -421 545 421
use sky130_fd_pr__pfet_01v8_8WDS2C  XM2
timestamp 1754378775
transform 1 0 2149 0 1 -123
box -545 -421 545 421
use sky130_fd_pr__pfet_01v8_8WDS2C  XM3
timestamp 1754378775
transform 1 0 2149 0 1 -859
box -545 -421 545 421
use sky130_fd_pr__pfet_01v8_8WDS2C  XM4
timestamp 1754378775
transform 1 0 1165 0 1 -1595
box -545 -421 545 421
use sky130_fd_pr__pfet_01v8_8WDS2C  XM5
timestamp 1754378775
transform 1 0 2149 0 1 -1595
box -545 -421 545 421
use sky130_fd_pr__pfet_01v8_8WDS2C  XM17
timestamp 1754378775
transform 1 0 1165 0 1 -123
box -545 -421 545 421
<< labels >>
flabel metal1 22 456 222 656 0 FreeSans 256 0 0 0 Vdd
port 1 nsew
flabel metal1 262 -2326 462 -2126 0 FreeSans 256 0 0 0 Vss
port 3 nsew
flabel metal1 2758 -590 2958 -390 0 FreeSans 256 0 0 0 Vref1
port 2 nsew
flabel metal1 2754 -1118 2952 -918 0 FreeSans 256 0 0 0 Vref2
port 0 nsew
flabel metal1 2768 -1376 2968 -1176 0 FreeSans 256 0 0 0 Vref3
port 4 nsew
flabel metal1 2740 -1848 2940 -1648 0 FreeSans 256 0 0 0 Vref4
port 5 nsew
rlabel metal1 948 -136 964 -106 1 lmid
<< end >>
