magic
tech sky130A
timestamp 1755358163
<< viali >>
rect 602 268 622 287
rect 602 60 631 83
<< metal1 >>
rect 412 537 512 637
rect 639 564 739 664
rect 439 432 470 537
rect 432 420 470 432
rect 432 402 463 420
rect 323 186 361 399
rect 423 360 428 402
rect 470 393 475 402
rect 470 371 557 393
rect 470 360 475 371
rect 645 370 669 564
rect 745 402 776 433
rect 731 360 736 402
rect 778 360 783 402
rect 432 325 463 360
rect 745 326 776 360
rect 595 287 640 291
rect 595 268 602 287
rect 622 271 640 287
rect 622 268 638 271
rect 438 222 469 229
rect 595 226 638 268
rect 437 188 471 222
rect 593 211 639 226
rect 595 196 639 211
rect 411 187 471 188
rect 407 186 436 187
rect 323 158 436 186
rect 323 150 361 158
rect 407 157 436 158
rect 471 157 476 187
rect 594 185 639 196
rect 738 194 769 225
rect 551 160 677 185
rect 437 131 471 157
rect 594 149 639 160
rect 732 156 737 194
rect 777 156 782 194
rect 438 122 469 131
rect 595 110 639 149
rect 738 118 769 156
rect 857 154 888 390
rect 596 83 637 110
rect 596 60 602 83
rect 631 60 637 83
rect 596 3 637 60
rect 571 -75 670 3
rect 570 -97 670 -75
<< via1 >>
rect 428 360 470 402
rect 736 360 778 402
rect 436 157 471 187
rect 737 156 777 194
<< metal2 >>
rect 428 402 470 407
rect 736 402 778 407
rect 470 361 736 384
rect 428 355 470 360
rect 778 361 779 384
rect 736 355 778 360
rect 737 194 777 199
rect 436 187 471 192
rect 430 160 436 187
rect 471 186 519 187
rect 471 185 546 186
rect 690 185 737 186
rect 471 161 737 185
rect 471 160 519 161
rect 690 157 737 161
rect 436 152 471 157
rect 737 151 777 156
use sky130_fd_pr__nfet_01v8_FEQNLY  XM1
timestamp 1754378775
transform 1 0 458 0 1 380
box -178 -130 178 130
use sky130_fd_pr__nfet_01v8_FEQNLY  XM2
timestamp 1754378775
transform 1 0 761 0 1 380
box -178 -130 178 130
use sky130_fd_pr__nfet_01v8_FEQNLY  XM3
timestamp 1754378775
transform 1 0 458 0 1 173
box -178 -130 178 130
use sky130_fd_pr__nfet_01v8_FEQNLY  XM4
timestamp 1754378775
transform 1 0 761 0 1 173
box -178 -130 178 130
<< labels >>
flabel metal1 412 537 512 637 0 FreeSans 128 0 0 0 Iin
port 0 nsew
flabel metal1 639 564 739 664 0 FreeSans 128 0 0 0 Iout
port 1 nsew
flabel metal1 571 -97 670 3 0 FreeSans 128 0 0 0 Vss
port 2 nsew
<< end >>
