magic
tech sky130A
magscale 1 2
timestamp 1755359579
<< locali >>
rect 858 -4748 3324 -4712
rect 858 -4826 954 -4748
rect 3238 -4826 3324 -4748
rect 858 -4856 3324 -4826
rect 3528 -4738 5508 -4716
rect 3528 -4842 3624 -4738
rect 5354 -4842 5508 -4738
rect 3528 -4866 5508 -4842
<< viali >>
rect 1976 472 2040 514
rect 1980 40 2032 74
rect 954 -4826 3238 -4748
rect 3624 -4842 5354 -4738
<< metal1 >>
rect 1932 1198 2132 1230
rect 1650 1042 2338 1198
rect 1656 348 1720 1042
rect 1932 1030 2132 1042
rect 1924 606 2124 806
rect 1962 514 2052 606
rect 1962 472 1976 514
rect 2040 472 2052 514
rect 1398 246 1530 286
rect 1018 74 1218 122
rect 1398 74 1430 246
rect 1668 172 1706 348
rect 1962 294 2052 472
rect 2266 324 2330 1042
rect 1882 260 2116 294
rect 1018 -20 1430 74
rect 1018 -78 1218 -20
rect 1398 -274 1430 -20
rect 1482 134 1714 172
rect 1482 -184 1512 134
rect 1966 74 2052 260
rect 2280 146 2318 324
rect 2504 272 2646 276
rect 2492 246 2646 272
rect 2504 244 2646 246
rect 2376 136 2540 168
rect 1966 40 1980 74
rect 2032 40 2052 74
rect 1966 18 2052 40
rect 1664 -274 1702 -54
rect 1398 -282 1702 -274
rect 1398 -302 1670 -282
rect 1428 -692 1628 -630
rect 1892 -692 1954 -146
rect 1428 -806 1954 -692
rect 1428 -830 1628 -806
rect 1794 -1718 1856 -1490
rect 1892 -1732 1954 -806
rect 2080 -666 2120 -122
rect 2278 -272 2316 -44
rect 2500 -188 2536 136
rect 2596 -6 2646 244
rect 2768 -6 2968 56
rect 2596 -100 2968 -6
rect 2596 -260 2646 -100
rect 2768 -144 2968 -100
rect 2446 -290 2646 -260
rect 2446 -292 2610 -290
rect 2328 -666 2528 -604
rect 2080 -780 2528 -666
rect 2080 -1066 2120 -780
rect 2328 -804 2528 -780
rect 2730 -1066 4170 -1058
rect 4466 -1066 4544 -1060
rect 2080 -1128 4544 -1066
rect 2182 -1132 4544 -1128
rect 2730 -1138 4170 -1132
rect 4466 -1618 4544 -1132
rect 2932 -4296 4912 -3972
rect 3170 -4708 3406 -4296
rect 3170 -4710 3522 -4708
rect 866 -4714 4680 -4710
rect 866 -4738 5508 -4714
rect 866 -4748 3624 -4738
rect 866 -4826 954 -4748
rect 3238 -4826 3624 -4748
rect 866 -4842 3624 -4826
rect 5354 -4842 5508 -4738
rect 866 -4848 5508 -4842
rect 3170 -4858 5508 -4848
rect 3322 -4866 5508 -4858
rect 3322 -4870 4382 -4866
rect 3322 -4908 3522 -4870
use sky130_fd_pr__res_generic_po_F4UD2D  R1
timestamp 1754378775
transform 1 0 4472 0 1 -2904
box -1166 -1596 1166 1596
use sky130_fd_pr__res_generic_po_F4UD2D  R2
timestamp 1754378775
transform 1 0 2118 0 1 -2918
box -1166 -1596 1166 1596
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM5
timestamp 1754378775
transform 1 0 1702 0 1 269
box -356 -269 356 269
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM6
timestamp 1754378775
transform 1 0 2308 0 1 -163
box -356 -269 356 269
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM7
timestamp 1754378775
transform 1 0 2308 0 1 269
box -356 -269 356 269
use sky130_fd_pr__pfet_01v8_CQSSBJ  XM11
timestamp 1754378775
transform 1 0 1702 0 1 -163
box -356 -269 356 269
<< labels >>
flabel metal1 1924 606 2124 806 0 FreeSans 256 0 0 0 Vdd
port 0 nsew
flabel metal1 3322 -4908 3522 -4708 0 FreeSans 256 0 0 0 Vss
port 1 nsew
flabel metal1 1932 1030 2132 1230 0 FreeSans 256 0 0 0 Ibias
port 6 nsew
flabel metal1 1428 -830 1628 -630 0 FreeSans 256 0 0 0 Iout1
port 2 nsew
flabel metal1 2328 -804 2528 -604 0 FreeSans 256 0 0 0 Iout2
port 3 nsew
flabel metal1 1018 -78 1218 122 0 FreeSans 256 0 0 0 Iin1
port 4 nsew
flabel metal1 2768 -144 2968 56 0 FreeSans 256 0 0 0 Iin2
port 5 nsew
<< end >>
