magic
tech sky130A
magscale 1 2
timestamp 1756317880
<< metal1 >>
rect 18186 42952 18196 42990
rect 17834 42906 18196 42952
rect 17828 42872 18196 42906
rect 17828 42444 17964 42872
rect 18186 42824 18196 42872
rect 18352 42952 18362 42990
rect 18352 42872 19144 42952
rect 18352 42824 18362 42872
rect 15834 42320 17964 42444
rect 17828 42314 17964 42320
rect 7926 41530 14058 41554
rect 7820 41524 14058 41530
rect 7820 41414 14398 41524
rect 7820 41400 14058 41414
rect 7820 38854 8438 41400
rect 16838 41192 17038 41244
rect 16838 41190 16888 41192
rect 16242 41070 16888 41190
rect 16838 41068 16888 41070
rect 16994 41068 17038 41192
rect 16838 41044 17038 41068
rect 15576 40326 15680 40846
rect 29406 40718 29680 40752
rect 21572 40686 29680 40718
rect 20992 40576 29680 40686
rect 21562 40538 29680 40576
rect 21572 40534 21628 40538
rect 21962 40534 29680 40538
rect 15464 39952 15474 40326
rect 15806 40184 15816 40326
rect 15806 40088 18602 40184
rect 15806 39952 15816 40088
rect 7756 38276 8438 38854
rect 29256 39682 29680 40534
rect 7756 37418 8430 38276
rect 9318 37484 9328 38012
rect 9954 37484 9964 38012
rect 7756 37290 8438 37418
rect 7820 35162 8438 37290
rect 7820 34108 8456 35162
rect 7824 33718 8456 34108
rect 11112 33942 11286 34726
rect 14810 33756 14984 34682
rect 19290 33834 19482 34702
rect 7820 33288 8456 33718
rect 10822 33430 10832 33598
rect 10964 33430 10974 33598
rect 11066 33596 11266 33616
rect 11066 33450 11080 33596
rect 11220 33450 11266 33596
rect 12272 33456 12390 33606
rect 18562 33570 18762 33592
rect 20456 33590 21112 33594
rect 11066 33416 11266 33450
rect 7824 32898 8456 33288
rect 7820 32834 8456 32898
rect 12270 33288 12390 33456
rect 13938 33482 14138 33506
rect 16828 33502 16954 33510
rect 13938 33320 13956 33482
rect 14110 33452 14138 33482
rect 14110 33360 14698 33452
rect 15948 33438 16954 33502
rect 15948 33410 16958 33438
rect 14110 33320 14138 33360
rect 13938 33306 14138 33320
rect 7820 30562 8438 32834
rect 12270 32766 12388 33288
rect 12270 32518 12390 32766
rect 16826 32656 16958 33410
rect 18562 33436 18610 33570
rect 18760 33528 18770 33570
rect 18760 33438 19142 33528
rect 20456 33506 21212 33590
rect 18760 33436 18770 33438
rect 18562 33392 18762 33436
rect 19054 33040 19284 33124
rect 12272 32282 12390 32518
rect 16828 32512 16954 32656
rect 21088 32556 21212 33506
rect 23714 31910 23866 33100
rect 23998 32132 24732 32174
rect 22442 31860 23866 31910
rect 22426 31818 23866 31860
rect 23994 32078 24732 32132
rect 22426 31808 23854 31818
rect 22426 31378 22578 31808
rect 23994 31612 24074 32078
rect 22416 31306 22578 31378
rect 23988 31550 24074 31612
rect 22416 31254 22534 31306
rect 21690 30974 21890 30992
rect 23988 30988 24062 31550
rect 21690 30968 22324 30974
rect 21690 30804 21726 30968
rect 21878 30832 22324 30968
rect 23584 30900 24062 30988
rect 23584 30888 23942 30900
rect 21878 30804 21890 30832
rect 21690 30792 21890 30804
rect 7820 30356 8430 30562
rect 22290 30454 22394 30530
rect 7798 28642 8430 30356
rect 22264 29596 22420 30454
rect 26070 30192 26080 30610
rect 26340 30192 26350 30610
rect 7820 27608 8430 28642
rect 12070 28494 14280 28508
rect 12038 28478 14280 28494
rect 18628 28478 18638 28510
rect 12038 28086 18638 28478
rect 12038 28022 14280 28086
rect 7820 20020 8438 27608
rect 11326 20400 11336 20980
rect 11750 20566 11760 20980
rect 12038 20566 12510 28022
rect 18628 27990 18638 28086
rect 18996 27990 19006 28510
rect 26080 28288 26304 30192
rect 29256 28502 29642 39682
rect 29256 28356 29638 28502
rect 26024 28216 26034 28288
rect 26010 28054 26034 28216
rect 26024 27906 26034 28054
rect 26392 27906 26402 28288
rect 26066 27486 26362 27906
rect 27286 27572 29654 28356
rect 19090 27242 26362 27486
rect 19102 25154 19240 27242
rect 26066 27208 26362 27242
rect 19108 24510 19234 25154
rect 19108 24388 19238 24510
rect 12916 22748 12926 22934
rect 13078 22748 13088 22934
rect 19126 21434 19238 24388
rect 19504 22782 19514 22934
rect 19660 22782 19670 22934
rect 17756 21292 19240 21434
rect 14596 20822 14606 20938
rect 14732 20822 14742 20938
rect 11750 20562 12898 20566
rect 11750 20446 13728 20562
rect 16620 20516 16820 20518
rect 16620 20500 17496 20516
rect 16620 20480 17512 20500
rect 11750 20400 11760 20446
rect 12038 20432 13728 20446
rect 15444 20422 17512 20480
rect 16620 20338 17512 20422
rect 16620 20318 16820 20338
rect 7822 19722 8438 20020
rect 7822 19718 11892 19722
rect 12500 19718 12510 19744
rect 7822 19620 12510 19718
rect 7784 19590 11892 19620
rect 7784 19562 8438 19590
rect 12500 19568 12510 19620
rect 12704 19568 12714 19744
rect 7784 10214 8238 19562
rect 12556 18646 12566 18876
rect 12918 18646 12928 18876
rect 11818 18534 12016 18540
rect 15810 18534 15820 18610
rect 11818 18356 15820 18534
rect 11818 14022 12016 18356
rect 15810 18342 15820 18356
rect 16046 18342 16056 18610
rect 13030 17088 13040 17250
rect 13232 17088 13242 17250
rect 14536 15152 14546 15282
rect 14676 15152 14686 15282
rect 12238 14724 12248 14902
rect 12402 14866 12412 14902
rect 12402 14736 13594 14866
rect 17378 14854 17512 20338
rect 17756 19476 17910 21292
rect 17732 19208 17910 19476
rect 18262 20962 18492 20976
rect 18816 20962 18826 21060
rect 18262 20890 18826 20962
rect 17732 17402 17886 19208
rect 12402 14724 12412 14736
rect 15422 14726 17512 14854
rect 17378 14702 17512 14726
rect 17720 17252 17886 17402
rect 17720 15370 17874 17252
rect 11804 13960 12576 14022
rect 15412 13994 15500 14394
rect 15410 13882 15500 13994
rect 17720 14036 17888 15370
rect 18262 15100 18492 20890
rect 18816 20850 18826 20890
rect 19006 20850 19016 21060
rect 19126 20664 19238 21292
rect 21174 20850 21184 20994
rect 21296 20850 21306 20994
rect 27328 20988 27850 27572
rect 19158 20592 19238 20664
rect 19158 20454 20246 20592
rect 27328 20150 27786 20988
rect 21964 20052 27786 20150
rect 27328 20006 27786 20052
rect 19052 19612 19062 19744
rect 19218 19612 19228 19744
rect 19088 18690 19098 18920
rect 19450 18690 19460 18920
rect 23622 17782 23822 17812
rect 19126 17596 19136 17738
rect 19284 17596 19294 17738
rect 22350 17612 23822 17782
rect 22350 17602 23742 17612
rect 20880 15646 20890 15772
rect 21006 15646 21016 15772
rect 19846 15212 19856 15370
rect 20014 15212 20024 15370
rect 27346 15362 27764 20006
rect 21772 15176 27786 15362
rect 18296 14562 18492 15100
rect 18296 14432 19044 14562
rect 18296 14412 18492 14432
rect 15410 13562 15498 13882
rect 17720 13836 18596 14036
rect 18704 13836 18746 14036
rect 17720 13810 18746 13836
rect 15352 13400 15362 13562
rect 15520 13400 15530 13562
rect 12556 12982 12566 13186
rect 12758 12982 12768 13186
rect 18908 13126 19082 13628
rect 16834 13016 19082 13126
rect 16834 12998 18876 13016
rect 18286 12710 18410 12756
rect 17076 12620 17086 12668
rect 14620 12482 17086 12620
rect 14622 12110 14752 12482
rect 17076 12388 17086 12482
rect 17384 12388 17394 12668
rect 18196 12480 18206 12710
rect 18484 12480 18494 12710
rect 18286 12366 18410 12480
rect 17518 12274 18410 12366
rect 17512 12214 18410 12274
rect 15096 12118 15774 12204
rect 7784 10076 8226 10214
rect 7758 9910 8226 10076
rect 7720 9848 8226 9910
rect 7720 9456 7784 9848
rect 8200 9456 8226 9848
rect 7720 9418 8226 9456
rect 14888 4992 15094 10924
rect 15656 10618 15768 12118
rect 17512 11884 17644 12214
rect 18286 12202 18410 12214
rect 17970 11858 18728 12010
rect 15656 10544 15780 10618
rect 15668 8312 15780 10544
rect 17838 10306 17936 10634
rect 17604 9934 17614 10306
rect 18018 9934 18028 10306
rect 16512 9292 16522 9518
rect 16762 9292 16772 9518
rect 16516 8878 16526 9074
rect 16734 8878 16744 9074
rect 18526 8308 18728 11858
rect 20516 9972 20526 10326
rect 20796 10268 20806 10326
rect 20796 9972 20818 10268
rect 17402 8144 18728 8308
rect 15466 7598 15666 7640
rect 15466 7488 15504 7598
rect 15620 7564 15666 7598
rect 17530 7608 17730 7658
rect 17530 7584 17556 7608
rect 15620 7488 16146 7564
rect 16994 7530 17556 7584
rect 15466 7470 16146 7488
rect 17530 7498 17556 7530
rect 17672 7498 17730 7608
rect 15466 7440 15666 7470
rect 17530 7458 17730 7498
rect 14342 3336 14352 3658
rect 14750 3520 14760 3658
rect 14902 3542 15094 4992
rect 20636 3560 20818 9972
rect 14902 3520 17108 3542
rect 14750 3402 17108 3520
rect 14750 3336 14760 3402
rect 14902 3400 17108 3402
rect 20058 3396 20818 3560
<< via1 >>
rect 18196 42824 18352 42990
rect 16888 41068 16994 41192
rect 15474 39952 15806 40326
rect 9328 37484 9954 38012
rect 10832 33430 10964 33598
rect 11080 33450 11220 33596
rect 13956 33320 14110 33482
rect 18610 33436 18760 33570
rect 21726 30804 21878 30968
rect 26080 30192 26340 30610
rect 11336 20400 11750 20980
rect 18638 27990 18996 28510
rect 26034 27906 26392 28288
rect 12926 22748 13078 22934
rect 19514 22782 19660 22934
rect 14606 20822 14732 20938
rect 12510 19568 12704 19744
rect 12566 18646 12918 18876
rect 15820 18342 16046 18610
rect 13040 17088 13232 17250
rect 14546 15152 14676 15282
rect 12248 14724 12402 14902
rect 18826 20850 19006 21060
rect 21184 20850 21296 20994
rect 19062 19612 19218 19744
rect 19098 18690 19450 18920
rect 19136 17596 19284 17738
rect 20890 15646 21006 15772
rect 19856 15212 20014 15370
rect 18596 13836 18704 14036
rect 15362 13400 15520 13562
rect 12566 12982 12758 13186
rect 17086 12388 17384 12668
rect 18206 12480 18484 12710
rect 7784 9456 8200 9848
rect 17614 9934 18018 10306
rect 16522 9292 16762 9518
rect 16526 8878 16734 9074
rect 20526 9972 20796 10326
rect 15504 7488 15620 7598
rect 17556 7498 17672 7608
rect 14352 3336 14750 3658
<< metal2 >>
rect 22372 43652 29418 43674
rect 16880 43610 29418 43652
rect 16880 43600 29440 43610
rect 16880 43440 29218 43600
rect 16880 43430 29440 43440
rect 16880 43422 29418 43430
rect 16888 41202 16986 43422
rect 22372 43420 29418 43422
rect 18196 42990 18352 43000
rect 18196 42814 18352 42824
rect 16888 41192 16994 41202
rect 16888 41058 16994 41068
rect 15474 40326 15806 40336
rect 15474 39942 15806 39952
rect 9328 38012 9954 38022
rect 9328 37474 9954 37484
rect 10832 33598 10964 33608
rect 10824 33588 10832 33598
rect 10964 33588 10966 33598
rect 11080 33596 11220 33606
rect 18610 33570 18760 33580
rect 11080 33440 11220 33450
rect 13956 33482 14110 33492
rect 10824 33418 10966 33428
rect 18610 33426 18760 33436
rect 13956 33310 14110 33320
rect 21726 30968 21878 30978
rect 21726 30794 21878 30804
rect 26080 30610 26340 30620
rect 26080 30182 26340 30192
rect 18594 28520 18978 29094
rect 18594 28510 18996 28520
rect 18594 28400 18638 28510
rect 18588 28094 18638 28400
rect 18638 27980 18996 27990
rect 26034 28288 26392 28298
rect 26034 27896 26392 27906
rect 12926 22934 13078 22944
rect 19514 22934 19660 22944
rect 19514 22772 19660 22782
rect 12926 22738 13078 22748
rect 18826 21060 19006 21070
rect 11336 20980 11750 20990
rect 14606 20938 14732 20948
rect 15880 20906 15982 20912
rect 14732 20822 15982 20906
rect 21184 20994 21296 21004
rect 19006 20886 21184 20958
rect 18826 20840 19006 20850
rect 21184 20840 21296 20850
rect 14606 20812 14732 20822
rect 11336 20390 11750 20400
rect 15880 20736 15982 20822
rect 11502 14830 11632 20390
rect 15880 20074 15984 20736
rect 12510 19744 12704 19754
rect 12510 19558 12704 19568
rect 12566 18876 12918 18886
rect 12566 18636 12918 18646
rect 15876 18868 15984 20074
rect 19062 19744 19218 19754
rect 19062 19602 19218 19612
rect 19098 18920 19450 18930
rect 15876 18620 15980 18868
rect 19098 18680 19450 18690
rect 15820 18610 16046 18620
rect 15820 18332 16046 18342
rect 19136 17738 19284 17748
rect 19136 17586 19284 17596
rect 13040 17250 13232 17260
rect 13040 17078 13232 17088
rect 20890 15772 21006 15782
rect 18246 15646 20890 15756
rect 18246 15636 21006 15646
rect 18246 15604 18708 15636
rect 18278 15544 18438 15604
rect 17114 15292 17338 15308
rect 14546 15282 17348 15292
rect 14676 15152 17348 15282
rect 14546 15142 14676 15152
rect 12248 14902 12402 14912
rect 11502 14748 12248 14830
rect 12402 14748 12436 14830
rect 12248 14714 12402 14724
rect 15362 13562 15520 13572
rect 15362 13390 15520 13400
rect 12534 13206 12794 13216
rect 12534 12968 12794 12978
rect 17114 12678 17338 15152
rect 18260 14412 18438 15544
rect 19856 15370 20014 15380
rect 18588 15212 19856 15354
rect 18588 15202 20014 15212
rect 18588 15186 19990 15202
rect 18260 13470 18418 14412
rect 18596 14036 18738 15186
rect 18704 13836 18738 14036
rect 18596 13826 18704 13836
rect 18260 13324 18438 13470
rect 18278 12720 18438 13324
rect 18206 12710 18484 12720
rect 17086 12668 17384 12678
rect 18206 12470 18484 12480
rect 17086 12378 17384 12388
rect 20526 10326 20796 10336
rect 17614 10306 18018 10316
rect 18018 10042 20526 10256
rect 20526 9962 20796 9972
rect 17614 9924 18018 9934
rect 7784 9848 8200 9858
rect 8200 9582 11366 9596
rect 8200 9528 16750 9582
rect 8200 9518 16762 9528
rect 8200 9456 16522 9518
rect 7784 9446 16522 9456
rect 7810 9418 16522 9446
rect 7910 9406 11366 9418
rect 16522 9282 16762 9292
rect 16526 9074 16734 9084
rect 16526 8868 16734 8878
rect 12568 7630 12888 7644
rect 22528 7638 22694 7642
rect 21988 7632 22850 7638
rect 21988 7630 22528 7632
rect 12568 7608 15608 7630
rect 17542 7608 22528 7630
rect 12568 7598 15620 7608
rect 12568 7488 15504 7598
rect 17542 7520 17556 7608
rect 17672 7520 22528 7608
rect 21928 7510 22528 7520
rect 22694 7510 22850 7632
rect 21928 7504 22850 7510
rect 21928 7498 22156 7504
rect 22528 7500 22694 7504
rect 17556 7488 17672 7498
rect 12568 7478 15620 7488
rect 12568 7432 15608 7478
rect 12568 2526 12888 7432
rect 14352 3658 14750 3668
rect 14352 3326 14750 3336
rect 25190 2526 25576 2536
rect 12542 2242 25190 2526
rect 12542 2232 25576 2242
rect 12542 2208 25486 2232
<< via2 >>
rect 29218 43440 29440 43600
rect 18196 42824 18352 42990
rect 15474 39952 15806 40326
rect 9328 37484 9954 38012
rect 10824 33430 10832 33588
rect 10832 33430 10964 33588
rect 10964 33430 10966 33588
rect 11080 33450 11220 33596
rect 10824 33428 10966 33430
rect 13956 33320 14110 33482
rect 18610 33436 18760 33570
rect 21726 30804 21878 30968
rect 12926 22748 13078 22934
rect 19514 22782 19660 22934
rect 12510 19568 12704 19744
rect 12566 18646 12918 18876
rect 19062 19612 19218 19744
rect 19098 18690 19450 18920
rect 19136 17596 19284 17738
rect 13040 17088 13232 17250
rect 15362 13400 15520 13562
rect 12534 13186 12794 13206
rect 12534 12982 12566 13186
rect 12566 12982 12758 13186
rect 12758 12982 12794 13186
rect 12534 12978 12794 12982
rect 16526 8878 16734 9074
rect 22528 7510 22694 7632
rect 14352 3336 14750 3658
rect 25190 2242 25576 2526
<< metal3 >>
rect 29166 43800 29176 44044
rect 29472 43800 29482 44044
rect 29218 43605 29428 43800
rect 29208 43600 29450 43605
rect 29208 43440 29218 43600
rect 29440 43440 29450 43600
rect 29208 43435 29450 43440
rect 18186 42990 18362 42995
rect 18186 42824 18196 42990
rect 18352 42824 18362 42990
rect 18186 42819 18362 42824
rect 23962 42428 24286 42436
rect 23946 42042 23956 42428
rect 24270 42042 24286 42428
rect 4414 40212 4424 40354
rect 4354 40048 4424 40212
rect 4414 39924 4424 40048
rect 4752 40212 4762 40354
rect 15464 40326 15816 40331
rect 6516 40212 6914 40250
rect 4752 40210 7124 40212
rect 15464 40210 15474 40326
rect 4752 40114 15474 40210
rect 4752 40048 7124 40114
rect 4752 39924 4762 40048
rect 15464 39952 15474 40114
rect 15806 40210 15816 40326
rect 15806 40114 16224 40210
rect 15806 39952 15816 40114
rect 15464 39947 15816 39952
rect 23962 39142 24286 42042
rect 24720 42012 24730 42398
rect 25044 42012 25054 42398
rect 11306 39128 24314 39142
rect 10804 38936 24314 39128
rect 10804 38892 12090 38936
rect 9318 38012 9964 38017
rect 9318 37484 9328 38012
rect 9954 37484 9964 38012
rect 9318 37479 9964 37484
rect 10804 33593 10968 38892
rect 13992 38748 14168 38778
rect 13964 38734 17274 38748
rect 24810 38734 24974 42012
rect 25378 41942 25388 42328
rect 25702 41942 25712 42328
rect 25792 41956 25802 42342
rect 26116 41956 26126 42342
rect 13964 38542 25010 38734
rect 11070 33596 11230 33601
rect 10804 33588 10976 33593
rect 10804 33428 10824 33588
rect 10966 33582 10976 33588
rect 11070 33582 11080 33596
rect 10966 33450 11080 33582
rect 11220 33450 11230 33596
rect 13992 33487 14168 38542
rect 15942 38514 25010 38542
rect 24810 38496 24974 38514
rect 18622 38420 18782 38436
rect 18622 38376 19090 38420
rect 25478 38384 25602 41942
rect 25838 40384 26060 41956
rect 21768 38376 25602 38384
rect 18622 38260 25602 38376
rect 18622 33575 18782 38260
rect 21768 38250 25602 38260
rect 21758 38096 21902 38112
rect 25780 38096 26114 40384
rect 21744 37822 26142 38096
rect 10966 33445 11230 33450
rect 13946 33482 14168 33487
rect 10966 33432 11210 33445
rect 10966 33428 10976 33432
rect 10804 33423 10976 33428
rect 10804 33398 10968 33423
rect 13946 33320 13956 33482
rect 14110 33320 14168 33482
rect 18600 33570 18782 33575
rect 18600 33436 18610 33570
rect 18760 33476 18782 33570
rect 18760 33436 18770 33476
rect 18600 33431 18770 33436
rect 13946 33315 14168 33320
rect 13992 33298 14168 33315
rect 21758 30973 21902 37822
rect 21716 30968 21902 30973
rect 21716 30804 21726 30968
rect 21878 30804 21902 30968
rect 21716 30799 21888 30804
rect 12916 22934 13088 22939
rect 12916 22748 12926 22934
rect 13078 22748 13088 22934
rect 19504 22934 19670 22939
rect 19504 22782 19514 22934
rect 19660 22782 19670 22934
rect 19504 22777 19670 22782
rect 12916 22743 13088 22748
rect 12500 19744 12714 19749
rect 12500 19568 12510 19744
rect 12704 19730 12714 19744
rect 19052 19744 19228 19749
rect 19052 19730 19062 19744
rect 12704 19612 19062 19730
rect 19218 19612 19228 19744
rect 12704 19607 19228 19612
rect 12704 19568 19224 19607
rect 12500 19563 12714 19568
rect 4380 18646 4390 18930
rect 4794 18892 7198 18930
rect 19088 18920 19460 18925
rect 19088 18892 19098 18920
rect 4794 18876 19098 18892
rect 4794 18672 12566 18876
rect 4794 18646 7198 18672
rect 12556 18646 12566 18672
rect 12918 18690 19098 18876
rect 19450 18892 19460 18920
rect 19450 18690 24096 18892
rect 12918 18672 24096 18690
rect 12918 18646 12928 18672
rect 12556 18641 12928 18646
rect 19126 17738 19294 17743
rect 19126 17596 19136 17738
rect 19284 17596 19294 17738
rect 19126 17591 19294 17596
rect 13040 17255 13050 17256
rect 13030 17250 13050 17255
rect 13030 17088 13040 17250
rect 13242 17094 13252 17256
rect 13232 17088 13242 17094
rect 13030 17083 13242 17088
rect 15352 13562 15530 13567
rect 15352 13542 15362 13562
rect 15284 13400 15362 13542
rect 15520 13542 15530 13562
rect 29328 13542 30550 13590
rect 15520 13400 30550 13542
rect 15284 13308 30550 13400
rect 29328 13292 30550 13308
rect 12466 13206 12808 13214
rect 4380 12606 4390 13000
rect 4826 12950 4836 13000
rect 12466 12978 12534 13206
rect 12794 12978 12808 13206
rect 6516 12958 8956 12966
rect 12466 12958 12808 12978
rect 6516 12950 12808 12958
rect 4826 12828 12808 12950
rect 4826 12606 12818 12828
rect 6516 12602 12818 12606
rect 16516 9074 16744 9079
rect 16516 8878 16526 9074
rect 16734 8878 16744 9074
rect 16516 8873 16744 8878
rect 22518 7634 22704 7637
rect 22516 7632 22712 7634
rect 22516 7510 22528 7632
rect 22694 7510 22712 7632
rect 22516 7308 22712 7510
rect 6516 3814 6586 3920
rect 4198 3806 6586 3814
rect 7976 3806 15316 3858
rect 4198 3742 15316 3806
rect 4198 3334 4340 3742
rect 4330 3300 4340 3334
rect 4678 3658 15316 3742
rect 4678 3336 14352 3658
rect 14750 3336 15316 3658
rect 4678 3334 15316 3336
rect 4678 3300 4688 3334
rect 6516 3320 15316 3334
rect 6516 3316 7928 3320
rect 22512 2162 22722 7308
rect 25180 2526 25586 2531
rect 26416 2526 26426 2548
rect 25180 2242 25190 2526
rect 25576 2242 26426 2526
rect 25180 2237 25586 2242
rect 26416 2208 26426 2242
rect 26744 2208 26754 2548
rect 22426 1720 22436 2162
rect 22900 1720 22910 2162
rect 30304 2096 30536 13292
rect 30282 1756 30292 2096
rect 30610 1756 30620 2096
<< via3 >>
rect 29176 43800 29472 44044
rect 18196 42824 18352 42990
rect 23956 42042 24270 42428
rect 4424 39924 4752 40354
rect 24730 42012 25044 42398
rect 9328 37484 9954 38012
rect 25388 41942 25702 42328
rect 25802 41956 26116 42342
rect 12926 22748 13078 22934
rect 19514 22782 19660 22934
rect 4390 18646 4794 18930
rect 19136 17596 19284 17738
rect 13050 17250 13242 17256
rect 13050 17094 13232 17250
rect 13232 17094 13242 17250
rect 4390 12606 4826 13000
rect 16526 8878 16734 9074
rect 4340 3300 4678 3742
rect 26426 2208 26744 2548
rect 22436 1720 22900 2162
rect 30292 1756 30610 2096
<< metal4 >>
rect 6132 44952 6194 45152
rect 6686 44952 6746 45152
rect 7236 44952 7298 45152
rect 7790 44952 7850 45152
rect 8340 44952 8402 45152
rect 8894 45150 8954 45152
rect 8892 44950 8954 45150
rect 9446 44952 9506 45152
rect 9924 44992 9984 45158
rect 9916 44902 9998 44992
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19996 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 45024 26066 45152
rect 26558 45038 26620 45152
rect 26004 44718 26066 45024
rect 26552 44952 26620 45038
rect 27108 45012 27170 45152
rect 27660 45080 27722 45152
rect 27108 44952 27176 45012
rect 26552 44738 26614 44952
rect 27114 44872 27176 44952
rect 23968 44560 26066 44718
rect 23968 44556 25926 44560
rect 4410 40354 4810 43932
rect 4410 39924 4424 40354
rect 4752 39924 4810 40354
rect 4410 18931 4810 39924
rect 5302 42976 5702 43946
rect 6292 42976 6998 42994
rect 18195 42990 18353 42991
rect 5302 42970 7394 42976
rect 10006 42970 11552 42982
rect 18195 42970 18196 42990
rect 5302 42824 18196 42970
rect 18352 42970 18353 42990
rect 18352 42824 19124 42970
rect 5302 42770 19124 42824
rect 5302 42732 7394 42770
rect 10006 42766 11552 42770
rect 5302 38276 5702 42732
rect 6292 42718 6998 42732
rect 23968 42429 24216 44556
rect 24802 44316 24950 44322
rect 26550 44316 26616 44738
rect 24802 44312 26618 44316
rect 24802 44156 26630 44312
rect 24802 44154 26618 44156
rect 23955 42428 24271 42429
rect 23955 42042 23956 42428
rect 24270 42042 24271 42428
rect 24802 42399 24950 44154
rect 27098 44036 27176 44872
rect 27650 44952 27722 45080
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 45068 29378 45152
rect 29310 44964 29394 45068
rect 27650 44820 27712 44952
rect 27650 44730 27722 44820
rect 27656 44476 27722 44730
rect 25894 44034 27180 44036
rect 25452 43932 27180 44034
rect 25452 43906 26088 43932
rect 23955 42041 24271 42042
rect 24729 42398 25045 42399
rect 24729 42012 24730 42398
rect 25044 42012 25045 42398
rect 25466 42329 25614 43906
rect 26070 43788 27548 43792
rect 27634 43788 27734 44476
rect 29284 44045 29412 44964
rect 29175 44044 29473 44045
rect 29175 43800 29176 44044
rect 29472 43800 29473 44044
rect 29175 43799 29473 43800
rect 26070 43772 27734 43788
rect 25882 43662 27734 43772
rect 25882 43660 27322 43662
rect 25882 42343 26008 43660
rect 25801 42342 26117 42343
rect 24729 42011 25045 42012
rect 25387 42328 25703 42329
rect 25387 41942 25388 42328
rect 25702 41942 25703 42328
rect 25801 41956 25802 42342
rect 26116 41956 26117 42342
rect 25801 41955 26117 41956
rect 25387 41941 25703 41942
rect 5302 37916 5678 38276
rect 9327 38012 9955 38013
rect 9327 37916 9328 38012
rect 5302 37898 9328 37916
rect 5282 37508 9328 37898
rect 5282 37500 5678 37508
rect 4389 18930 4810 18931
rect 4389 18646 4390 18930
rect 4794 18646 4810 18930
rect 4389 18645 4810 18646
rect 4410 13001 4810 18645
rect 5302 37418 5678 37500
rect 9327 37484 9328 37508
rect 9954 37916 9955 38012
rect 9954 37508 10002 37916
rect 9954 37484 9955 37508
rect 9327 37483 9955 37484
rect 5302 34108 5702 37418
rect 5302 33718 5656 34108
rect 5302 22960 5702 33718
rect 6292 22960 7110 23020
rect 5302 22908 7110 22960
rect 12925 22934 13079 22935
rect 12925 22908 12926 22934
rect 5302 22756 12926 22908
rect 5302 22698 7110 22756
rect 12925 22748 12926 22756
rect 13078 22908 13079 22934
rect 19513 22934 19661 22935
rect 19513 22908 19514 22934
rect 13078 22796 19514 22908
rect 13078 22756 13168 22796
rect 19513 22782 19514 22796
rect 19660 22908 19661 22934
rect 19660 22796 19758 22908
rect 19660 22782 19661 22796
rect 19513 22781 19661 22782
rect 13078 22748 13079 22756
rect 12925 22747 13079 22748
rect 5302 17448 5702 22698
rect 6292 22642 7110 22698
rect 12984 17738 19986 17772
rect 12984 17610 19136 17738
rect 5274 17292 7718 17448
rect 13018 17292 13264 17610
rect 19135 17596 19136 17610
rect 19284 17610 19986 17738
rect 19284 17596 19285 17610
rect 19135 17595 19285 17596
rect 5274 17256 13318 17292
rect 5274 17094 13050 17256
rect 13242 17094 13318 17256
rect 5274 17034 13318 17094
rect 5274 16908 7718 17034
rect 4389 13000 4827 13001
rect 4389 12606 4390 13000
rect 4826 12606 4827 13000
rect 4389 12605 4827 12606
rect 4410 3743 4810 12605
rect 4339 3742 4810 3743
rect 4339 3300 4340 3742
rect 4678 3300 4810 3742
rect 4339 3299 4810 3300
rect 4410 780 4810 3299
rect 5302 9226 5702 16908
rect 5302 9090 8016 9226
rect 5302 9074 17076 9090
rect 5302 8878 16526 9074
rect 16734 8878 17076 9074
rect 5302 8768 17076 8878
rect 5302 8686 8016 8768
rect 5302 794 5702 8686
rect 26425 2548 26745 2549
rect 26425 2208 26426 2548
rect 26744 2208 26745 2548
rect 26425 2207 26745 2208
rect 22435 2162 22901 2163
rect 22435 1720 22436 2162
rect 22900 1720 22901 2162
rect 26472 1720 26664 2207
rect 30291 2096 30611 2097
rect 30291 1756 30292 2096
rect 30610 1756 30611 2096
rect 30291 1755 30611 1756
rect 22435 1719 22901 1720
rect 22656 200 22800 1719
rect 26512 200 26656 1720
rect 30382 204 30526 1755
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30360 194 30546 204
rect 30356 8 30546 194
rect 30356 -2 30542 8
use dac_tt  x1
timestamp 1755904430
transform 1 0 -2232 0 1 29998
box 11390 -1060 31196 7786
use bump_final_tt  x2
timestamp 1755119682
transform 1 0 11464 0 1 16782
box 986 -3802 5584 490
use vol_ref_gen_tt  x3
timestamp 1755355673
transform 1 0 18162 0 1 42354
box 22 -2326 2968 656
use ccm_nmos_tt  x4
timestamp 1755358163
transform 1 0 16640 0 1 10714
box 560 -194 1878 1328
use bump_final_tt  x5
timestamp 1755119682
transform 1 0 11520 0 1 22458
box 986 -3802 5584 490
use bump_final_tt  x6
timestamp 1755119682
transform 1 0 18064 0 1 22506
box 986 -3802 5584 490
use bump_final_tt  x7
timestamp 1755119682
transform 1 0 17794 0 1 17286
box 986 -3802 5584 490
use ccm_nmos_tt  x8
timestamp 1755358163
transform 1 0 13758 0 1 10946
box 560 -194 1878 1328
use inv_layout_tt  x9
timestamp 1755205548
transform 1 0 15584 0 1 34482
box -1072 -1780 500 -190
use inv_layout_tt  x10
timestamp 1755205548
transform 1 0 11882 0 1 34604
box -1072 -1780 500 -190
use ref_gen_tt  x11
timestamp 1755360409
transform 1 0 14450 0 1 41668
box -156 -944 1886 810
use wta_pmos_tt  x12
timestamp 1755359579
transform 1 0 14608 0 1 8268
box 858 -4908 5638 1230
use inv_layout_tt  x13
timestamp 1755205548
transform 1 0 20078 0 1 34588
box -1072 -1780 500 -190
use inv_layout_tt  x14
timestamp 1755205548
transform 1 0 23194 0 1 31992
box -1072 -1780 500 -190
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel via1 14456 3418 14656 3618 0 FreeSans 256 0 0 0 Vss
port 1 nsew
flabel metal1 16838 41044 17038 41244 0 FreeSans 256 0 0 0 En
port 7 nsew
flabel metal4 s 9924 44958 9984 45158 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal1 16620 20318 16820 20518 0 FreeSans 256 0 0 0 Vr
port 2 nsew
flabel metal1 15466 7440 15666 7640 0 FreeSans 256 0 0 0 Iout0
port 8 nsew
flabel metal1 17530 7458 17730 7658 0 FreeSans 256 0 0 0 Iout1
port 9 nsew
flabel metal1 23622 17612 23822 17812 0 FreeSans 256 0 0 0 Vdd
port 0 nsew
flabel metal4 5302 794 5656 43946 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 4410 780 4810 43932 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal1 21690 30792 21700 30992 0 FreeSans 256 0 0 0 Vin1
port 6 nsew
flabel metal1 18562 33392 18762 33592 0 FreeSans 256 0 0 0 Vin2
port 5 nsew
flabel metal1 13938 33306 14138 33506 0 FreeSans 256 0 0 0 Vin3
port 4 nsew
flabel metal1 11066 33416 11266 33616 0 FreeSans 256 0 0 0 Vin4
port 3 nsew
rlabel metal1 13318 41436 13430 41512 1 Ibias
rlabel metal1 29328 39956 29586 40310 1 Vref4
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
