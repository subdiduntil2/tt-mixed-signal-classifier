magic
tech sky130A
magscale 1 2
timestamp 1755120335
<< locali >>
rect 1096 418 2134 436
rect 1096 368 1216 418
rect 2112 368 2134 418
rect 1096 356 2134 368
<< viali >>
rect 1216 368 2112 418
rect 1594 228 1632 262
rect 1166 -966 1202 -932
rect 1958 -970 2000 -926
<< metal1 >>
rect 958 436 1158 456
rect 958 418 2134 436
rect 958 384 1216 418
rect 632 368 1216 384
rect 2112 412 2134 418
rect 2112 410 2214 412
rect 2112 380 2294 410
rect 2112 368 2134 380
rect 632 356 2134 368
rect 632 306 1158 356
rect 632 -528 708 306
rect 958 256 1158 306
rect 1560 288 1652 356
rect 1562 262 1652 288
rect 1562 228 1594 262
rect 1632 238 1652 262
rect 1632 228 1654 238
rect 1562 200 1654 228
rect 1502 156 1674 164
rect 1814 156 1862 164
rect 1502 120 1862 156
rect 1502 114 1674 120
rect 934 -76 1134 26
rect 1194 -76 1204 -34
rect 934 -112 1204 -76
rect 934 -174 1134 -112
rect 1194 -128 1204 -112
rect 1268 -128 1278 -34
rect 1544 -126 1554 -24
rect 1640 -126 1650 -24
rect 1814 -106 1862 120
rect 1958 -106 2158 -52
rect 1814 -154 2158 -106
rect 1428 -230 1438 -196
rect 1424 -314 1438 -230
rect 1498 -314 1508 -196
rect 1670 -310 1680 -192
rect 1740 -310 1750 -192
rect 632 -562 1212 -528
rect 632 -592 1214 -562
rect 484 -716 684 -646
rect 484 -780 774 -716
rect 484 -846 684 -780
rect 764 -786 774 -780
rect 830 -786 840 -716
rect 1150 -888 1214 -592
rect 1424 -662 1468 -314
rect 1814 -472 1862 -154
rect 1958 -252 2158 -154
rect 2232 -398 2292 380
rect 2232 -440 2290 -398
rect 1506 -508 1862 -472
rect 1506 -522 1678 -508
rect 1814 -510 1862 -508
rect 1944 -502 2290 -440
rect 1422 -700 1574 -662
rect 1472 -702 1574 -700
rect 1134 -932 1214 -888
rect 1134 -966 1166 -932
rect 1202 -966 1214 -932
rect 1134 -978 1214 -966
rect 1544 -802 1574 -702
rect 720 -1044 1290 -1040
rect 720 -1072 1398 -1044
rect 720 -1076 1290 -1072
rect 720 -1278 756 -1076
rect 648 -1478 848 -1278
rect 1262 -1312 1272 -1186
rect 1374 -1312 1384 -1186
rect 704 -1664 764 -1478
rect 1156 -1526 1166 -1438
rect 1238 -1526 1248 -1438
rect 1394 -1522 1404 -1434
rect 1476 -1480 1486 -1434
rect 1544 -1480 1572 -802
rect 1944 -926 2028 -502
rect 2514 -784 2714 -698
rect 2160 -846 2170 -786
rect 2236 -848 2714 -784
rect 2514 -898 2714 -848
rect 1944 -970 1958 -926
rect 2000 -970 2028 -926
rect 1944 -980 2028 -970
rect 2376 -1038 2428 -1036
rect 1818 -1046 2428 -1038
rect 1720 -1074 2428 -1046
rect 1818 -1080 2428 -1074
rect 1738 -1302 1748 -1208
rect 1826 -1302 1836 -1208
rect 2376 -1316 2428 -1080
rect 1622 -1480 1632 -1420
rect 1476 -1516 1632 -1480
rect 1476 -1522 1486 -1516
rect 1622 -1530 1632 -1516
rect 1704 -1530 1714 -1420
rect 1856 -1530 1866 -1420
rect 1938 -1530 1948 -1420
rect 2278 -1516 2478 -1316
rect 2362 -1662 2398 -1516
rect 704 -1670 1280 -1664
rect 704 -1680 1392 -1670
rect 1840 -1676 2398 -1662
rect 704 -1698 1398 -1680
rect 704 -1708 1280 -1698
rect 1724 -1704 2398 -1676
rect 884 -1710 1280 -1708
<< via1 >>
rect 1204 -128 1268 -34
rect 1554 -126 1640 -24
rect 1438 -314 1498 -196
rect 1680 -310 1740 -192
rect 774 -786 830 -716
rect 1272 -1312 1374 -1186
rect 1166 -1526 1238 -1438
rect 1404 -1522 1476 -1434
rect 2170 -846 2236 -786
rect 1748 -1302 1826 -1208
rect 1632 -1530 1704 -1420
rect 1866 -1530 1938 -1420
<< metal2 >>
rect 1554 -24 1640 -14
rect 1204 -34 1268 -24
rect 1268 -110 1554 -56
rect 1204 -138 1268 -128
rect 1554 -136 1640 -126
rect 1438 -196 1498 -186
rect 1680 -192 1740 -182
rect 1498 -286 1680 -238
rect 1438 -324 1498 -314
rect 1680 -320 1740 -310
rect 774 -716 830 -706
rect 830 -726 1342 -716
rect 830 -784 1344 -726
rect 774 -796 830 -786
rect 1300 -1176 1344 -784
rect 2170 -786 2236 -776
rect 1760 -844 2170 -786
rect 1272 -1186 1374 -1176
rect 1762 -1198 1802 -844
rect 2170 -856 2236 -846
rect 1748 -1208 1826 -1198
rect 1748 -1312 1826 -1302
rect 1272 -1322 1374 -1312
rect 1632 -1420 1704 -1410
rect 1166 -1438 1238 -1428
rect 1404 -1434 1476 -1424
rect 1238 -1506 1404 -1458
rect 1166 -1536 1238 -1526
rect 1404 -1532 1476 -1522
rect 1866 -1420 1938 -1410
rect 1704 -1504 1866 -1452
rect 1632 -1540 1704 -1530
rect 1866 -1540 1938 -1530
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM3
timestamp 1754378775
transform 1 0 1319 0 1 -1375
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM5
timestamp 1754378775
transform 1 0 1783 0 1 -1375
box -285 -469 285 469
use sky130_fd_pr__pfet_01v8_JMP7WZ  XM8
timestamp 1754378775
transform 1 0 1587 0 1 -179
box -285 -469 285 469
<< labels >>
flabel metal1 648 -1478 848 -1278 0 FreeSans 256 0 0 0 Vin
port 3 nsew
flabel metal1 2278 -1516 2478 -1316 0 FreeSans 256 0 0 0 Vindot
port 4 nsew
flabel metal1 1958 -252 2158 -52 0 FreeSans 256 0 0 0 Vg
port 1 nsew
flabel metal1 2514 -898 2714 -698 0 FreeSans 256 0 0 0 Vout2
port 6 nsew
flabel metal1 484 -846 684 -646 0 FreeSans 256 0 0 0 Vout1
port 5 nsew
flabel metal1 934 -174 1134 26 0 FreeSans 256 0 0 0 Vupper
port 0 nsew
flabel metal1 958 256 1158 456 0 FreeSans 256 0 0 0 Vdd
port 2 nsew
rlabel metal1 1492 -696 1534 -670 1 l1
<< end >>
